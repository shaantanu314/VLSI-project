magic
tech scmos
timestamp 1618572623
<< ntransistor >>
rect -3 109 -1 119
rect -33 98 -31 108
rect -94 87 -92 97
rect -57 88 -55 98
rect 58 95 60 105
rect -33 73 -31 83
rect 58 70 60 80
rect 34 38 36 48
rect -121 11 -119 21
<< ptransistor >>
rect -94 111 -92 131
rect -33 120 -31 140
rect 58 117 60 137
rect -57 54 -55 74
rect -3 75 -1 95
rect 34 62 36 82
rect -121 33 -119 53
rect -33 41 -31 61
rect 58 38 60 58
<< ndiffusion >>
rect -4 109 -3 119
rect -1 109 0 119
rect -34 98 -33 108
rect -31 98 -30 108
rect -95 87 -94 97
rect -92 87 -91 97
rect -58 88 -57 98
rect -55 88 -54 98
rect 57 95 58 105
rect 60 95 61 105
rect -34 73 -33 83
rect -31 73 -30 83
rect 57 70 58 80
rect 60 70 61 80
rect 33 38 34 48
rect 36 38 37 48
rect -122 11 -121 21
rect -119 11 -118 21
<< pdiffusion >>
rect -95 111 -94 131
rect -92 111 -91 131
rect -34 120 -33 140
rect -31 120 -30 140
rect 57 117 58 137
rect 60 117 61 137
rect -58 54 -57 74
rect -55 54 -54 74
rect -4 75 -3 95
rect -1 75 0 95
rect 33 62 34 82
rect 36 62 37 82
rect -122 33 -121 53
rect -119 33 -118 53
rect -34 41 -33 61
rect -31 41 -30 61
rect 57 38 58 58
rect 60 38 61 58
<< ndcontact >>
rect -8 109 -4 119
rect 0 109 4 119
rect -38 98 -34 108
rect -30 98 -26 108
rect -99 87 -95 97
rect -91 87 -87 97
rect -62 88 -58 98
rect -54 88 -50 98
rect 53 95 57 105
rect 61 95 65 105
rect -38 73 -34 83
rect -30 73 -26 83
rect 53 70 57 80
rect 61 70 65 80
rect 29 38 33 48
rect 37 38 41 48
rect -126 11 -122 21
rect -118 11 -114 21
<< pdcontact >>
rect -99 111 -95 131
rect -91 111 -87 131
rect -38 120 -34 140
rect -30 120 -26 140
rect 53 117 57 137
rect 61 117 65 137
rect -62 54 -58 74
rect -54 54 -50 74
rect -8 75 -4 95
rect 0 75 4 95
rect 29 62 33 82
rect 37 62 41 82
rect -126 33 -122 53
rect -118 33 -114 53
rect -38 41 -34 61
rect -30 41 -26 61
rect 53 38 57 58
rect 61 38 65 58
<< polysilicon >>
rect -33 140 -31 143
rect -94 131 -92 138
rect 58 137 60 140
rect -94 106 -92 111
rect -33 108 -31 120
rect -3 119 -1 126
rect -94 97 -92 102
rect -57 98 -55 105
rect -3 104 -1 109
rect 58 105 60 117
rect -33 95 -31 98
rect -3 95 -1 100
rect -94 80 -92 87
rect -57 83 -55 88
rect -33 83 -31 86
rect -57 74 -55 79
rect -121 53 -119 56
rect 58 92 60 95
rect 34 82 36 89
rect -33 61 -31 73
rect -3 68 -1 75
rect 58 80 60 83
rect -57 47 -55 54
rect 34 57 36 62
rect 58 58 60 70
rect 34 48 36 53
rect -33 38 -31 41
rect -121 21 -119 33
rect 34 31 36 38
rect 58 35 60 38
rect -121 8 -119 11
<< polycontact >>
rect -98 134 -94 138
rect -7 122 -3 126
rect -37 113 -33 117
rect 54 110 58 114
rect -61 101 -57 105
rect -98 80 -94 84
rect 30 85 34 89
rect -7 68 -3 72
rect -31 64 -27 68
rect -61 47 -57 51
rect 60 61 64 65
rect -125 26 -121 30
rect 30 31 34 35
<< metal1 >>
rect -41 145 -33 148
rect -38 140 -34 145
rect 50 142 58 145
rect -100 134 -98 138
rect -105 119 -99 123
rect -105 106 -102 119
rect -87 119 -81 123
rect 53 137 57 142
rect -10 122 -7 126
rect -113 103 -102 106
rect -105 94 -102 103
rect -84 106 -81 119
rect -30 117 -26 120
rect -75 113 -37 117
rect -30 113 -20 117
rect -75 106 -72 113
rect -30 108 -26 113
rect -84 103 -72 106
rect -105 90 -99 94
rect -84 94 -81 103
rect -87 90 -81 94
rect -105 80 -98 84
rect -129 58 -121 61
rect -126 53 -122 58
rect -131 26 -125 30
rect -118 29 -114 33
rect -105 51 -101 80
rect -75 71 -72 103
rect -63 101 -61 105
rect -23 103 -20 113
rect -14 112 -8 116
rect -14 103 -11 112
rect 4 112 10 116
rect 61 114 65 117
rect -23 100 -11 103
rect -68 91 -62 95
rect -68 71 -65 91
rect -50 91 -44 95
rect -75 68 -65 71
rect -68 66 -65 68
rect -68 62 -62 66
rect -47 68 -44 91
rect -38 92 -34 98
rect -38 89 -26 92
rect -30 83 -26 89
rect -38 68 -34 73
rect -23 69 -20 100
rect -14 87 -11 100
rect 7 96 10 112
rect 16 110 54 114
rect 61 110 71 114
rect 16 96 19 110
rect 61 105 65 110
rect -14 83 -8 87
rect 7 92 19 96
rect 7 87 10 92
rect 4 83 10 87
rect -24 68 -20 69
rect -47 66 -34 68
rect -50 64 -34 66
rect -27 64 -20 68
rect -14 68 -7 72
rect 16 68 19 92
rect 68 104 71 110
rect 68 101 76 104
rect 53 89 57 95
rect 27 85 30 89
rect 53 86 65 89
rect 23 70 29 74
rect 23 68 26 70
rect -50 62 -44 64
rect -38 61 -34 64
rect -105 47 -61 51
rect -105 29 -101 47
rect -30 36 -26 41
rect -31 33 -23 36
rect -14 35 -10 68
rect 16 65 26 68
rect 23 45 26 65
rect 61 80 65 86
rect 41 70 47 74
rect 44 65 47 70
rect 53 65 57 70
rect 68 66 71 101
rect 67 65 71 66
rect 44 61 57 65
rect 64 61 71 65
rect 23 41 29 45
rect 44 45 47 61
rect 41 41 47 45
rect 53 58 57 61
rect -14 31 30 35
rect 61 33 65 38
rect -14 29 -9 31
rect 60 30 68 33
rect -118 28 -113 29
rect -105 28 -9 29
rect -118 25 -9 28
rect -118 21 -114 25
rect -126 6 -122 11
<< labels >>
rlabel metal1 -128 28 -128 28 3 clk
rlabel metal1 -124 59 -124 59 1 vdd
rlabel metal1 -124 8 -124 8 1 gnd
rlabel metal1 -28 35 -28 35 1 vdd
rlabel metal1 -29 90 -29 90 1 gnd
rlabel metal1 -38 147 -38 147 5 vdd
rlabel metal1 -99 136 -99 136 1 clk
rlabel metal1 -62 102 -62 102 1 clk
rlabel metal1 53 144 53 144 5 vdd
rlabel metal1 62 87 62 87 1 gnd
rlabel metal1 63 32 63 32 1 vdd
rlabel metal1 28 87 28 87 3 clk
rlabel metal1 -9 123 -9 123 1 clk
rlabel metal1 -112 104 -112 104 1 D
rlabel metal1 74 102 74 102 7 Q
<< end >>
