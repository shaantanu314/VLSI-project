magic
tech scmos
timestamp 1619629090
<< error_p >>
rect -172 -762 -164 -761
<< ntransistor >>
rect 522 16 524 26
rect 492 5 494 15
rect 431 -6 433 4
rect 468 -5 470 5
rect 583 2 585 12
rect 492 -20 494 -10
rect 583 -23 585 -13
rect -132 -81 -130 -71
rect 559 -55 561 -45
rect -162 -92 -160 -82
rect 404 -82 406 -72
rect -223 -103 -221 -93
rect -186 -102 -184 -92
rect -71 -95 -69 -85
rect -162 -117 -160 -107
rect -71 -120 -69 -110
rect -95 -152 -93 -142
rect -250 -179 -248 -169
rect -133 -227 -131 -217
rect -163 -238 -161 -228
rect -224 -249 -222 -239
rect -187 -248 -185 -238
rect -72 -241 -70 -231
rect -163 -263 -161 -253
rect -3 -253 -1 -243
rect 11 -253 13 -243
rect 36 -244 38 -234
rect 50 -244 52 -234
rect -72 -266 -70 -256
rect 154 -246 156 -236
rect 168 -246 170 -236
rect 193 -237 195 -227
rect 207 -237 209 -227
rect 522 -244 524 -234
rect 76 -267 78 -257
rect 90 -267 92 -257
rect 233 -260 235 -250
rect 247 -260 249 -250
rect 492 -255 494 -245
rect -96 -298 -94 -288
rect 431 -266 433 -256
rect 468 -265 470 -255
rect 583 -258 585 -248
rect 36 -313 38 -303
rect 50 -313 52 -303
rect 193 -306 195 -296
rect 207 -306 209 -296
rect 492 -280 494 -270
rect 583 -283 585 -273
rect -251 -325 -249 -315
rect 559 -315 561 -305
rect -133 -368 -131 -358
rect 404 -342 406 -332
rect -163 -379 -161 -369
rect -224 -390 -222 -380
rect -187 -389 -185 -379
rect -72 -382 -70 -372
rect 29 -379 31 -369
rect 43 -379 45 -369
rect 63 -379 65 -369
rect -163 -404 -161 -394
rect -72 -407 -70 -397
rect 145 -403 147 -393
rect 159 -403 161 -393
rect 179 -403 181 -393
rect 219 -405 221 -395
rect 227 -405 229 -395
rect 244 -405 246 -395
rect -96 -439 -94 -429
rect -251 -466 -249 -456
rect -134 -511 -132 -501
rect -164 -522 -162 -512
rect -225 -533 -223 -523
rect -188 -532 -186 -522
rect -73 -525 -71 -515
rect -164 -547 -162 -537
rect 3 -538 5 -528
rect 17 -538 19 -528
rect 42 -529 44 -519
rect 56 -529 58 -519
rect -73 -550 -71 -540
rect 160 -531 162 -521
rect 174 -531 176 -521
rect 199 -522 201 -512
rect 213 -522 215 -512
rect 522 -528 524 -518
rect 82 -552 84 -542
rect 96 -552 98 -542
rect 239 -545 241 -535
rect 253 -545 255 -535
rect 492 -539 494 -529
rect -97 -582 -95 -572
rect 431 -550 433 -540
rect 468 -549 470 -539
rect 583 -542 585 -532
rect 42 -598 44 -588
rect 56 -598 58 -588
rect 199 -591 201 -581
rect 213 -591 215 -581
rect 492 -564 494 -554
rect 583 -567 585 -557
rect -252 -609 -250 -599
rect 559 -599 561 -589
rect -134 -652 -132 -642
rect 404 -626 406 -616
rect -164 -663 -162 -653
rect -225 -674 -223 -664
rect -188 -673 -186 -663
rect -73 -666 -71 -656
rect 35 -664 37 -654
rect 49 -664 51 -654
rect 69 -664 71 -654
rect -164 -688 -162 -678
rect -73 -691 -71 -681
rect 151 -688 153 -678
rect 165 -688 167 -678
rect 185 -688 187 -678
rect 224 -688 226 -678
rect 238 -688 240 -678
rect 258 -688 260 -678
rect 295 -690 297 -680
rect 303 -690 305 -680
rect 320 -690 322 -680
rect -97 -723 -95 -713
rect -252 -750 -250 -740
rect 248 -771 250 -761
rect 256 -771 258 -761
rect 273 -771 275 -761
rect -134 -800 -132 -790
rect -164 -811 -162 -801
rect 522 -797 524 -787
rect -225 -822 -223 -812
rect -188 -821 -186 -811
rect -73 -814 -71 -804
rect 492 -808 494 -798
rect -164 -836 -162 -826
rect 431 -819 433 -809
rect 468 -818 470 -808
rect 583 -811 585 -801
rect -73 -839 -71 -829
rect -97 -871 -95 -861
rect 492 -833 494 -823
rect 583 -836 585 -826
rect -252 -898 -250 -888
rect 559 -868 561 -858
rect -134 -941 -132 -931
rect 3 -918 5 -908
rect 17 -918 19 -908
rect 42 -909 44 -899
rect 56 -909 58 -899
rect 160 -911 162 -901
rect 174 -911 176 -901
rect 199 -902 201 -892
rect 213 -902 215 -892
rect 404 -895 406 -885
rect 82 -932 84 -922
rect 96 -932 98 -922
rect 239 -925 241 -915
rect 253 -925 255 -915
rect -164 -952 -162 -942
rect -225 -963 -223 -953
rect -188 -962 -186 -952
rect -73 -955 -71 -945
rect -164 -977 -162 -967
rect -73 -980 -71 -970
rect 42 -978 44 -968
rect 56 -978 58 -968
rect 199 -971 201 -961
rect 213 -971 215 -961
rect -97 -1012 -95 -1002
rect -252 -1039 -250 -1029
rect 35 -1044 37 -1034
rect 49 -1044 51 -1034
rect 69 -1044 71 -1034
rect 522 -1016 524 -1006
rect 492 -1027 494 -1017
rect 431 -1038 433 -1028
rect 468 -1037 470 -1027
rect 583 -1030 585 -1020
rect 151 -1068 153 -1058
rect 165 -1068 167 -1058
rect 185 -1068 187 -1058
rect 224 -1068 226 -1058
rect 238 -1068 240 -1058
rect 258 -1068 260 -1058
rect 296 -1070 298 -1060
rect 304 -1070 306 -1060
rect 321 -1070 323 -1060
rect 492 -1052 494 -1042
rect 583 -1055 585 -1045
rect 559 -1087 561 -1077
rect 404 -1114 406 -1104
rect 149 -1160 151 -1150
rect 163 -1160 165 -1150
rect 183 -1160 185 -1150
rect 215 -1162 217 -1152
rect 223 -1162 225 -1152
rect 240 -1162 242 -1152
rect 265 -1169 267 -1159
rect 273 -1169 275 -1159
rect 290 -1169 292 -1159
<< ptransistor >>
rect 431 18 433 38
rect 492 27 494 47
rect 583 24 585 44
rect 468 -39 470 -19
rect 522 -18 524 2
rect 559 -31 561 -11
rect -223 -79 -221 -59
rect -162 -70 -160 -50
rect -71 -73 -69 -53
rect 404 -60 406 -40
rect 492 -52 494 -32
rect 583 -55 585 -35
rect -186 -136 -184 -116
rect -132 -115 -130 -95
rect -95 -128 -93 -108
rect -250 -157 -248 -137
rect -162 -149 -160 -129
rect -71 -152 -69 -132
rect -224 -225 -222 -205
rect -163 -216 -161 -196
rect -72 -219 -70 -199
rect -3 -228 -1 -208
rect 11 -228 13 -208
rect 36 -219 38 -199
rect 50 -219 52 -199
rect -187 -282 -185 -262
rect -133 -261 -131 -241
rect 154 -221 156 -201
rect 168 -221 170 -201
rect 193 -212 195 -192
rect 207 -212 209 -192
rect 76 -242 78 -222
rect 90 -242 92 -222
rect -96 -274 -94 -254
rect 233 -235 235 -215
rect 247 -235 249 -215
rect 431 -242 433 -222
rect 492 -233 494 -213
rect 583 -236 585 -216
rect -251 -303 -249 -283
rect -163 -295 -161 -275
rect -72 -298 -70 -278
rect 36 -288 38 -268
rect 50 -288 52 -268
rect 193 -281 195 -261
rect 207 -281 209 -261
rect 468 -299 470 -279
rect 522 -278 524 -258
rect 559 -291 561 -271
rect 404 -320 406 -300
rect 492 -312 494 -292
rect 583 -315 585 -295
rect -224 -366 -222 -346
rect -163 -357 -161 -337
rect -72 -360 -70 -340
rect 29 -354 31 -334
rect 43 -354 45 -334
rect 63 -354 65 -334
rect 145 -378 147 -358
rect 159 -378 161 -358
rect 179 -378 181 -358
rect -187 -423 -185 -403
rect -133 -402 -131 -382
rect 219 -383 221 -363
rect 226 -383 228 -363
rect 244 -383 246 -363
rect -96 -415 -94 -395
rect -251 -444 -249 -424
rect -163 -436 -161 -416
rect -72 -439 -70 -419
rect -225 -509 -223 -489
rect -164 -500 -162 -480
rect -73 -503 -71 -483
rect 3 -513 5 -493
rect 17 -513 19 -493
rect 42 -504 44 -484
rect 56 -504 58 -484
rect -188 -566 -186 -546
rect -134 -545 -132 -525
rect 160 -506 162 -486
rect 174 -506 176 -486
rect 199 -497 201 -477
rect 213 -497 215 -477
rect -97 -558 -95 -538
rect 82 -527 84 -507
rect 96 -527 98 -507
rect 239 -520 241 -500
rect 253 -520 255 -500
rect 431 -526 433 -506
rect 492 -517 494 -497
rect 583 -520 585 -500
rect -252 -587 -250 -567
rect -164 -579 -162 -559
rect -73 -582 -71 -562
rect 42 -573 44 -553
rect 56 -573 58 -553
rect 199 -566 201 -546
rect 213 -566 215 -546
rect 468 -583 470 -563
rect 522 -562 524 -542
rect 559 -575 561 -555
rect 404 -604 406 -584
rect 492 -596 494 -576
rect 583 -599 585 -579
rect -225 -650 -223 -630
rect -164 -641 -162 -621
rect -73 -644 -71 -624
rect 35 -639 37 -619
rect 49 -639 51 -619
rect 69 -639 71 -619
rect 151 -663 153 -643
rect 165 -663 167 -643
rect 185 -663 187 -643
rect 224 -663 226 -643
rect 238 -663 240 -643
rect 258 -663 260 -643
rect -188 -707 -186 -687
rect -134 -686 -132 -666
rect 295 -668 297 -648
rect 302 -668 304 -648
rect 320 -668 322 -648
rect -97 -699 -95 -679
rect -252 -728 -250 -708
rect -164 -720 -162 -700
rect -73 -723 -71 -703
rect 248 -749 250 -729
rect 255 -749 257 -729
rect 273 -749 275 -729
rect -225 -798 -223 -778
rect -164 -789 -162 -769
rect -73 -792 -71 -772
rect 431 -795 433 -775
rect 492 -786 494 -766
rect 583 -789 585 -769
rect -188 -855 -186 -835
rect -134 -834 -132 -814
rect -97 -847 -95 -827
rect -252 -876 -250 -856
rect -164 -868 -162 -848
rect -73 -871 -71 -851
rect 468 -852 470 -832
rect 522 -831 524 -811
rect 559 -844 561 -824
rect 3 -893 5 -873
rect 17 -893 19 -873
rect 42 -884 44 -864
rect 56 -884 58 -864
rect 160 -886 162 -866
rect 174 -886 176 -866
rect 199 -877 201 -857
rect 213 -877 215 -857
rect 404 -873 406 -853
rect 492 -865 494 -845
rect 583 -868 585 -848
rect -225 -939 -223 -919
rect -164 -930 -162 -910
rect -73 -933 -71 -913
rect 82 -907 84 -887
rect 96 -907 98 -887
rect 239 -900 241 -880
rect 253 -900 255 -880
rect 42 -953 44 -933
rect 56 -953 58 -933
rect 199 -946 201 -926
rect 213 -946 215 -926
rect -188 -996 -186 -976
rect -134 -975 -132 -955
rect -97 -988 -95 -968
rect -252 -1017 -250 -997
rect -164 -1009 -162 -989
rect -73 -1012 -71 -992
rect 35 -1019 37 -999
rect 49 -1019 51 -999
rect 69 -1019 71 -999
rect 431 -1014 433 -994
rect 492 -1005 494 -985
rect 151 -1043 153 -1023
rect 165 -1043 167 -1023
rect 185 -1043 187 -1023
rect 224 -1043 226 -1023
rect 238 -1043 240 -1023
rect 258 -1043 260 -1023
rect 583 -1008 585 -988
rect 296 -1048 298 -1028
rect 303 -1048 305 -1028
rect 321 -1048 323 -1028
rect 468 -1071 470 -1051
rect 522 -1050 524 -1030
rect 559 -1063 561 -1043
rect 404 -1092 406 -1072
rect 492 -1084 494 -1064
rect 583 -1087 585 -1067
rect 149 -1135 151 -1115
rect 163 -1135 165 -1115
rect 183 -1135 185 -1115
rect 215 -1140 217 -1120
rect 222 -1140 224 -1120
rect 240 -1140 242 -1120
rect 265 -1147 267 -1127
rect 272 -1147 274 -1127
rect 290 -1147 292 -1127
<< ndiffusion >>
rect 521 16 522 26
rect 524 16 525 26
rect 491 5 492 15
rect 494 5 495 15
rect 430 -6 431 4
rect 433 -6 434 4
rect 467 -5 468 5
rect 470 -5 471 5
rect 582 2 583 12
rect 585 2 586 12
rect 491 -20 492 -10
rect 494 -20 495 -10
rect 582 -23 583 -13
rect 585 -23 586 -13
rect -133 -81 -132 -71
rect -130 -81 -129 -71
rect 558 -55 559 -45
rect 561 -55 562 -45
rect -163 -92 -162 -82
rect -160 -92 -159 -82
rect 403 -82 404 -72
rect 406 -82 407 -72
rect -224 -103 -223 -93
rect -221 -103 -220 -93
rect -187 -102 -186 -92
rect -184 -102 -183 -92
rect -72 -95 -71 -85
rect -69 -95 -68 -85
rect -163 -117 -162 -107
rect -160 -117 -159 -107
rect -72 -120 -71 -110
rect -69 -120 -68 -110
rect -96 -152 -95 -142
rect -93 -152 -92 -142
rect -251 -179 -250 -169
rect -248 -179 -247 -169
rect -134 -227 -133 -217
rect -131 -227 -130 -217
rect -164 -238 -163 -228
rect -161 -238 -160 -228
rect -225 -249 -224 -239
rect -222 -249 -221 -239
rect -188 -248 -187 -238
rect -185 -248 -184 -238
rect -73 -241 -72 -231
rect -70 -241 -69 -231
rect -164 -263 -163 -253
rect -161 -263 -160 -253
rect -4 -253 -3 -243
rect -1 -253 11 -243
rect 13 -253 14 -243
rect 35 -244 36 -234
rect 38 -244 50 -234
rect 52 -244 53 -234
rect -73 -266 -72 -256
rect -70 -266 -69 -256
rect 153 -246 154 -236
rect 156 -246 168 -236
rect 170 -246 171 -236
rect 192 -237 193 -227
rect 195 -237 207 -227
rect 209 -237 210 -227
rect 521 -244 522 -234
rect 524 -244 525 -234
rect 75 -267 76 -257
rect 78 -267 90 -257
rect 92 -267 93 -257
rect 232 -260 233 -250
rect 235 -260 247 -250
rect 249 -260 250 -250
rect 491 -255 492 -245
rect 494 -255 495 -245
rect -97 -298 -96 -288
rect -94 -298 -93 -288
rect 430 -266 431 -256
rect 433 -266 434 -256
rect 467 -265 468 -255
rect 470 -265 471 -255
rect 582 -258 583 -248
rect 585 -258 586 -248
rect 35 -313 36 -303
rect 38 -313 50 -303
rect 52 -313 53 -303
rect 192 -306 193 -296
rect 195 -306 207 -296
rect 209 -306 210 -296
rect 491 -280 492 -270
rect 494 -280 495 -270
rect 582 -283 583 -273
rect 585 -283 586 -273
rect -252 -325 -251 -315
rect -249 -325 -248 -315
rect 558 -315 559 -305
rect 561 -315 562 -305
rect -134 -368 -133 -358
rect -131 -368 -130 -358
rect 403 -342 404 -332
rect 406 -342 407 -332
rect -164 -379 -163 -369
rect -161 -379 -160 -369
rect -225 -390 -224 -380
rect -222 -390 -221 -380
rect -188 -389 -187 -379
rect -185 -389 -184 -379
rect -73 -382 -72 -372
rect -70 -382 -69 -372
rect 28 -379 29 -369
rect 31 -379 43 -369
rect 45 -379 46 -369
rect 60 -379 63 -369
rect 65 -379 68 -369
rect -164 -404 -163 -394
rect -161 -404 -160 -394
rect -73 -407 -72 -397
rect -70 -407 -69 -397
rect 144 -403 145 -393
rect 147 -403 159 -393
rect 161 -403 162 -393
rect 176 -403 179 -393
rect 181 -403 184 -393
rect 217 -405 219 -395
rect 221 -405 222 -395
rect 226 -405 227 -395
rect 229 -405 231 -395
rect 243 -405 244 -395
rect 246 -405 247 -395
rect -97 -439 -96 -429
rect -94 -439 -93 -429
rect -252 -466 -251 -456
rect -249 -466 -248 -456
rect -135 -511 -134 -501
rect -132 -511 -131 -501
rect -165 -522 -164 -512
rect -162 -522 -161 -512
rect -226 -533 -225 -523
rect -223 -533 -222 -523
rect -189 -532 -188 -522
rect -186 -532 -185 -522
rect -74 -525 -73 -515
rect -71 -525 -70 -515
rect -165 -547 -164 -537
rect -162 -547 -161 -537
rect 2 -538 3 -528
rect 5 -538 17 -528
rect 19 -538 20 -528
rect 41 -529 42 -519
rect 44 -529 56 -519
rect 58 -529 59 -519
rect -74 -550 -73 -540
rect -71 -550 -70 -540
rect 159 -531 160 -521
rect 162 -531 174 -521
rect 176 -531 177 -521
rect 198 -522 199 -512
rect 201 -522 213 -512
rect 215 -522 216 -512
rect 521 -528 522 -518
rect 524 -528 525 -518
rect 81 -552 82 -542
rect 84 -552 96 -542
rect 98 -552 99 -542
rect 238 -545 239 -535
rect 241 -545 253 -535
rect 255 -545 256 -535
rect 491 -539 492 -529
rect 494 -539 495 -529
rect -98 -582 -97 -572
rect -95 -582 -94 -572
rect 430 -550 431 -540
rect 433 -550 434 -540
rect 467 -549 468 -539
rect 470 -549 471 -539
rect 582 -542 583 -532
rect 585 -542 586 -532
rect 41 -598 42 -588
rect 44 -598 56 -588
rect 58 -598 59 -588
rect 198 -591 199 -581
rect 201 -591 213 -581
rect 215 -591 216 -581
rect 491 -564 492 -554
rect 494 -564 495 -554
rect 582 -567 583 -557
rect 585 -567 586 -557
rect -253 -609 -252 -599
rect -250 -609 -249 -599
rect 558 -599 559 -589
rect 561 -599 562 -589
rect -135 -652 -134 -642
rect -132 -652 -131 -642
rect 403 -626 404 -616
rect 406 -626 407 -616
rect -165 -663 -164 -653
rect -162 -663 -161 -653
rect -226 -674 -225 -664
rect -223 -674 -222 -664
rect -189 -673 -188 -663
rect -186 -673 -185 -663
rect -74 -666 -73 -656
rect -71 -666 -70 -656
rect 34 -664 35 -654
rect 37 -664 49 -654
rect 51 -664 52 -654
rect 66 -664 69 -654
rect 71 -664 74 -654
rect -165 -688 -164 -678
rect -162 -688 -161 -678
rect -74 -691 -73 -681
rect -71 -691 -70 -681
rect 150 -688 151 -678
rect 153 -688 165 -678
rect 167 -688 168 -678
rect 182 -688 185 -678
rect 187 -688 190 -678
rect 223 -688 224 -678
rect 226 -688 238 -678
rect 240 -688 241 -678
rect 255 -688 258 -678
rect 260 -688 263 -678
rect 293 -690 295 -680
rect 297 -690 298 -680
rect 302 -690 303 -680
rect 305 -690 307 -680
rect 319 -690 320 -680
rect 322 -690 323 -680
rect -98 -723 -97 -713
rect -95 -723 -94 -713
rect -253 -750 -252 -740
rect -250 -750 -249 -740
rect 246 -771 248 -761
rect 250 -771 251 -761
rect 255 -771 256 -761
rect 258 -771 260 -761
rect 272 -771 273 -761
rect 275 -771 276 -761
rect -135 -800 -134 -790
rect -132 -800 -131 -790
rect -165 -811 -164 -801
rect -162 -811 -161 -801
rect 521 -797 522 -787
rect 524 -797 525 -787
rect -226 -822 -225 -812
rect -223 -822 -222 -812
rect -189 -821 -188 -811
rect -186 -821 -185 -811
rect -74 -814 -73 -804
rect -71 -814 -70 -804
rect 491 -808 492 -798
rect 494 -808 495 -798
rect -165 -836 -164 -826
rect -162 -836 -161 -826
rect 430 -819 431 -809
rect 433 -819 434 -809
rect 467 -818 468 -808
rect 470 -818 471 -808
rect 582 -811 583 -801
rect 585 -811 586 -801
rect -74 -839 -73 -829
rect -71 -839 -70 -829
rect -98 -871 -97 -861
rect -95 -871 -94 -861
rect 491 -833 492 -823
rect 494 -833 495 -823
rect 582 -836 583 -826
rect 585 -836 586 -826
rect -253 -898 -252 -888
rect -250 -898 -249 -888
rect 558 -868 559 -858
rect 561 -868 562 -858
rect -135 -941 -134 -931
rect -132 -941 -131 -931
rect 2 -918 3 -908
rect 5 -918 17 -908
rect 19 -918 20 -908
rect 41 -909 42 -899
rect 44 -909 56 -899
rect 58 -909 59 -899
rect 159 -911 160 -901
rect 162 -911 174 -901
rect 176 -911 177 -901
rect 198 -902 199 -892
rect 201 -902 213 -892
rect 215 -902 216 -892
rect 403 -895 404 -885
rect 406 -895 407 -885
rect 81 -932 82 -922
rect 84 -932 96 -922
rect 98 -932 99 -922
rect 238 -925 239 -915
rect 241 -925 253 -915
rect 255 -925 256 -915
rect -165 -952 -164 -942
rect -162 -952 -161 -942
rect -226 -963 -225 -953
rect -223 -963 -222 -953
rect -189 -962 -188 -952
rect -186 -962 -185 -952
rect -74 -955 -73 -945
rect -71 -955 -70 -945
rect -165 -977 -164 -967
rect -162 -977 -161 -967
rect -74 -980 -73 -970
rect -71 -980 -70 -970
rect 41 -978 42 -968
rect 44 -978 56 -968
rect 58 -978 59 -968
rect 198 -971 199 -961
rect 201 -971 213 -961
rect 215 -971 216 -961
rect -98 -1012 -97 -1002
rect -95 -1012 -94 -1002
rect -253 -1039 -252 -1029
rect -250 -1039 -249 -1029
rect 34 -1044 35 -1034
rect 37 -1044 49 -1034
rect 51 -1044 52 -1034
rect 66 -1044 69 -1034
rect 71 -1044 74 -1034
rect 521 -1016 522 -1006
rect 524 -1016 525 -1006
rect 491 -1027 492 -1017
rect 494 -1027 495 -1017
rect 430 -1038 431 -1028
rect 433 -1038 434 -1028
rect 467 -1037 468 -1027
rect 470 -1037 471 -1027
rect 582 -1030 583 -1020
rect 585 -1030 586 -1020
rect 150 -1068 151 -1058
rect 153 -1068 165 -1058
rect 167 -1068 168 -1058
rect 182 -1068 185 -1058
rect 187 -1068 190 -1058
rect 223 -1068 224 -1058
rect 226 -1068 238 -1058
rect 240 -1068 241 -1058
rect 255 -1068 258 -1058
rect 260 -1068 263 -1058
rect 294 -1070 296 -1060
rect 298 -1070 299 -1060
rect 303 -1070 304 -1060
rect 306 -1070 308 -1060
rect 320 -1070 321 -1060
rect 323 -1070 324 -1060
rect 491 -1052 492 -1042
rect 494 -1052 495 -1042
rect 582 -1055 583 -1045
rect 585 -1055 586 -1045
rect 558 -1087 559 -1077
rect 561 -1087 562 -1077
rect 403 -1114 404 -1104
rect 406 -1114 407 -1104
rect 148 -1160 149 -1150
rect 151 -1160 163 -1150
rect 165 -1160 166 -1150
rect 180 -1160 183 -1150
rect 185 -1160 188 -1150
rect 213 -1162 215 -1152
rect 217 -1162 218 -1152
rect 222 -1162 223 -1152
rect 225 -1162 227 -1152
rect 239 -1162 240 -1152
rect 242 -1162 243 -1152
rect 263 -1169 265 -1159
rect 267 -1169 268 -1159
rect 272 -1169 273 -1159
rect 275 -1169 277 -1159
rect 289 -1169 290 -1159
rect 292 -1169 293 -1159
<< pdiffusion >>
rect 430 18 431 38
rect 433 18 434 38
rect 491 27 492 47
rect 494 27 495 47
rect 582 24 583 44
rect 585 24 586 44
rect 467 -39 468 -19
rect 470 -39 471 -19
rect 521 -18 522 2
rect 524 -18 525 2
rect 558 -31 559 -11
rect 561 -31 562 -11
rect -224 -79 -223 -59
rect -221 -79 -220 -59
rect -163 -70 -162 -50
rect -160 -70 -159 -50
rect -72 -73 -71 -53
rect -69 -73 -68 -53
rect 403 -60 404 -40
rect 406 -60 407 -40
rect 491 -52 492 -32
rect 494 -52 495 -32
rect 582 -55 583 -35
rect 585 -55 586 -35
rect -187 -136 -186 -116
rect -184 -136 -183 -116
rect -133 -115 -132 -95
rect -130 -115 -129 -95
rect -96 -128 -95 -108
rect -93 -128 -92 -108
rect -251 -157 -250 -137
rect -248 -157 -247 -137
rect -163 -149 -162 -129
rect -160 -149 -159 -129
rect -72 -152 -71 -132
rect -69 -152 -68 -132
rect -225 -225 -224 -205
rect -222 -225 -221 -205
rect -164 -216 -163 -196
rect -161 -216 -160 -196
rect -73 -219 -72 -199
rect -70 -219 -69 -199
rect -4 -228 -3 -208
rect -1 -228 3 -208
rect 7 -228 11 -208
rect 13 -228 14 -208
rect 35 -219 36 -199
rect 38 -219 42 -199
rect 46 -219 50 -199
rect 52 -219 53 -199
rect -188 -282 -187 -262
rect -185 -282 -184 -262
rect -134 -261 -133 -241
rect -131 -261 -130 -241
rect 153 -221 154 -201
rect 156 -221 160 -201
rect 164 -221 168 -201
rect 170 -221 171 -201
rect 192 -212 193 -192
rect 195 -212 199 -192
rect 203 -212 207 -192
rect 209 -212 210 -192
rect 75 -242 76 -222
rect 78 -242 82 -222
rect 86 -242 90 -222
rect 92 -242 93 -222
rect -97 -274 -96 -254
rect -94 -274 -93 -254
rect 232 -235 233 -215
rect 235 -235 239 -215
rect 243 -235 247 -215
rect 249 -235 250 -215
rect 430 -242 431 -222
rect 433 -242 434 -222
rect 491 -233 492 -213
rect 494 -233 495 -213
rect 582 -236 583 -216
rect 585 -236 586 -216
rect -252 -303 -251 -283
rect -249 -303 -248 -283
rect -164 -295 -163 -275
rect -161 -295 -160 -275
rect -73 -298 -72 -278
rect -70 -298 -69 -278
rect 35 -288 36 -268
rect 38 -288 42 -268
rect 46 -288 50 -268
rect 52 -288 53 -268
rect 192 -281 193 -261
rect 195 -281 199 -261
rect 203 -281 207 -261
rect 209 -281 210 -261
rect 467 -299 468 -279
rect 470 -299 471 -279
rect 521 -278 522 -258
rect 524 -278 525 -258
rect 558 -291 559 -271
rect 561 -291 562 -271
rect 403 -320 404 -300
rect 406 -320 407 -300
rect 491 -312 492 -292
rect 494 -312 495 -292
rect 582 -315 583 -295
rect 585 -315 586 -295
rect -225 -366 -224 -346
rect -222 -366 -221 -346
rect -164 -357 -163 -337
rect -161 -357 -160 -337
rect -73 -360 -72 -340
rect -70 -360 -69 -340
rect 28 -354 29 -334
rect 31 -354 35 -334
rect 39 -354 43 -334
rect 45 -354 46 -334
rect 60 -354 63 -334
rect 65 -354 68 -334
rect 144 -378 145 -358
rect 147 -378 151 -358
rect 155 -378 159 -358
rect 161 -378 162 -358
rect 176 -378 179 -358
rect 181 -378 184 -358
rect -188 -423 -187 -403
rect -185 -423 -184 -403
rect -134 -402 -133 -382
rect -131 -402 -130 -382
rect 217 -383 219 -363
rect 221 -383 226 -363
rect 228 -383 230 -363
rect 243 -383 244 -363
rect 246 -383 247 -363
rect -97 -415 -96 -395
rect -94 -415 -93 -395
rect -252 -444 -251 -424
rect -249 -444 -248 -424
rect -164 -436 -163 -416
rect -161 -436 -160 -416
rect -73 -439 -72 -419
rect -70 -439 -69 -419
rect -226 -509 -225 -489
rect -223 -509 -222 -489
rect -165 -500 -164 -480
rect -162 -500 -161 -480
rect -74 -503 -73 -483
rect -71 -503 -70 -483
rect 2 -513 3 -493
rect 5 -513 9 -493
rect 13 -513 17 -493
rect 19 -513 20 -493
rect 41 -504 42 -484
rect 44 -504 48 -484
rect 52 -504 56 -484
rect 58 -504 59 -484
rect -189 -566 -188 -546
rect -186 -566 -185 -546
rect -135 -545 -134 -525
rect -132 -545 -131 -525
rect 159 -506 160 -486
rect 162 -506 166 -486
rect 170 -506 174 -486
rect 176 -506 177 -486
rect 198 -497 199 -477
rect 201 -497 205 -477
rect 209 -497 213 -477
rect 215 -497 216 -477
rect -98 -558 -97 -538
rect -95 -558 -94 -538
rect 81 -527 82 -507
rect 84 -527 88 -507
rect 92 -527 96 -507
rect 98 -527 99 -507
rect 238 -520 239 -500
rect 241 -520 245 -500
rect 249 -520 253 -500
rect 255 -520 256 -500
rect 430 -526 431 -506
rect 433 -526 434 -506
rect 491 -517 492 -497
rect 494 -517 495 -497
rect 582 -520 583 -500
rect 585 -520 586 -500
rect -253 -587 -252 -567
rect -250 -587 -249 -567
rect -165 -579 -164 -559
rect -162 -579 -161 -559
rect -74 -582 -73 -562
rect -71 -582 -70 -562
rect 41 -573 42 -553
rect 44 -573 48 -553
rect 52 -573 56 -553
rect 58 -573 59 -553
rect 198 -566 199 -546
rect 201 -566 205 -546
rect 209 -566 213 -546
rect 215 -566 216 -546
rect 467 -583 468 -563
rect 470 -583 471 -563
rect 521 -562 522 -542
rect 524 -562 525 -542
rect 558 -575 559 -555
rect 561 -575 562 -555
rect 403 -604 404 -584
rect 406 -604 407 -584
rect 491 -596 492 -576
rect 494 -596 495 -576
rect 582 -599 583 -579
rect 585 -599 586 -579
rect -226 -650 -225 -630
rect -223 -650 -222 -630
rect -165 -641 -164 -621
rect -162 -641 -161 -621
rect -74 -644 -73 -624
rect -71 -644 -70 -624
rect 34 -639 35 -619
rect 37 -639 41 -619
rect 45 -639 49 -619
rect 51 -639 52 -619
rect 66 -639 69 -619
rect 71 -639 74 -619
rect 150 -663 151 -643
rect 153 -663 157 -643
rect 161 -663 165 -643
rect 167 -663 168 -643
rect 182 -663 185 -643
rect 187 -663 190 -643
rect 223 -663 224 -643
rect 226 -663 230 -643
rect 234 -663 238 -643
rect 240 -663 241 -643
rect 255 -663 258 -643
rect 260 -663 263 -643
rect -189 -707 -188 -687
rect -186 -707 -185 -687
rect -135 -686 -134 -666
rect -132 -686 -131 -666
rect 293 -668 295 -648
rect 297 -668 302 -648
rect 304 -668 306 -648
rect 319 -668 320 -648
rect 322 -668 323 -648
rect -98 -699 -97 -679
rect -95 -699 -94 -679
rect -253 -728 -252 -708
rect -250 -728 -249 -708
rect -165 -720 -164 -700
rect -162 -720 -161 -700
rect -74 -723 -73 -703
rect -71 -723 -70 -703
rect 246 -749 248 -729
rect 250 -749 255 -729
rect 257 -749 259 -729
rect 272 -749 273 -729
rect 275 -749 276 -729
rect -226 -798 -225 -778
rect -223 -798 -222 -778
rect -165 -789 -164 -769
rect -162 -789 -161 -769
rect -74 -792 -73 -772
rect -71 -792 -70 -772
rect 430 -795 431 -775
rect 433 -795 434 -775
rect 491 -786 492 -766
rect 494 -786 495 -766
rect 582 -789 583 -769
rect 585 -789 586 -769
rect -189 -855 -188 -835
rect -186 -855 -185 -835
rect -135 -834 -134 -814
rect -132 -834 -131 -814
rect -98 -847 -97 -827
rect -95 -847 -94 -827
rect -253 -876 -252 -856
rect -250 -876 -249 -856
rect -165 -868 -164 -848
rect -162 -868 -161 -848
rect -74 -871 -73 -851
rect -71 -871 -70 -851
rect 467 -852 468 -832
rect 470 -852 471 -832
rect 521 -831 522 -811
rect 524 -831 525 -811
rect 558 -844 559 -824
rect 561 -844 562 -824
rect 2 -893 3 -873
rect 5 -893 9 -873
rect 13 -893 17 -873
rect 19 -893 20 -873
rect 41 -884 42 -864
rect 44 -884 48 -864
rect 52 -884 56 -864
rect 58 -884 59 -864
rect 159 -886 160 -866
rect 162 -886 166 -866
rect 170 -886 174 -866
rect 176 -886 177 -866
rect 198 -877 199 -857
rect 201 -877 205 -857
rect 209 -877 213 -857
rect 215 -877 216 -857
rect 403 -873 404 -853
rect 406 -873 407 -853
rect 491 -865 492 -845
rect 494 -865 495 -845
rect 582 -868 583 -848
rect 585 -868 586 -848
rect -226 -939 -225 -919
rect -223 -939 -222 -919
rect -165 -930 -164 -910
rect -162 -930 -161 -910
rect -74 -933 -73 -913
rect -71 -933 -70 -913
rect 81 -907 82 -887
rect 84 -907 88 -887
rect 92 -907 96 -887
rect 98 -907 99 -887
rect 238 -900 239 -880
rect 241 -900 245 -880
rect 249 -900 253 -880
rect 255 -900 256 -880
rect 41 -953 42 -933
rect 44 -953 48 -933
rect 52 -953 56 -933
rect 58 -953 59 -933
rect 198 -946 199 -926
rect 201 -946 205 -926
rect 209 -946 213 -926
rect 215 -946 216 -926
rect -189 -996 -188 -976
rect -186 -996 -185 -976
rect -135 -975 -134 -955
rect -132 -975 -131 -955
rect -98 -988 -97 -968
rect -95 -988 -94 -968
rect -253 -1017 -252 -997
rect -250 -1017 -249 -997
rect -165 -1009 -164 -989
rect -162 -1009 -161 -989
rect -74 -1012 -73 -992
rect -71 -1012 -70 -992
rect 34 -1019 35 -999
rect 37 -1019 41 -999
rect 45 -1019 49 -999
rect 51 -1019 52 -999
rect 66 -1019 69 -999
rect 71 -1019 74 -999
rect 430 -1014 431 -994
rect 433 -1014 434 -994
rect 491 -1005 492 -985
rect 494 -1005 495 -985
rect 150 -1043 151 -1023
rect 153 -1043 157 -1023
rect 161 -1043 165 -1023
rect 167 -1043 168 -1023
rect 182 -1043 185 -1023
rect 187 -1043 190 -1023
rect 223 -1043 224 -1023
rect 226 -1043 230 -1023
rect 234 -1043 238 -1023
rect 240 -1043 241 -1023
rect 255 -1043 258 -1023
rect 260 -1043 263 -1023
rect 582 -1008 583 -988
rect 585 -1008 586 -988
rect 294 -1048 296 -1028
rect 298 -1048 303 -1028
rect 305 -1048 307 -1028
rect 320 -1048 321 -1028
rect 323 -1048 324 -1028
rect 467 -1071 468 -1051
rect 470 -1071 471 -1051
rect 521 -1050 522 -1030
rect 524 -1050 525 -1030
rect 558 -1063 559 -1043
rect 561 -1063 562 -1043
rect 403 -1092 404 -1072
rect 406 -1092 407 -1072
rect 491 -1084 492 -1064
rect 494 -1084 495 -1064
rect 582 -1087 583 -1067
rect 585 -1087 586 -1067
rect 148 -1135 149 -1115
rect 151 -1135 155 -1115
rect 159 -1135 163 -1115
rect 165 -1135 166 -1115
rect 180 -1135 183 -1115
rect 185 -1135 188 -1115
rect 213 -1140 215 -1120
rect 217 -1140 222 -1120
rect 224 -1140 226 -1120
rect 239 -1140 240 -1120
rect 242 -1140 243 -1120
rect 263 -1147 265 -1127
rect 267 -1147 272 -1127
rect 274 -1147 276 -1127
rect 289 -1147 290 -1127
rect 292 -1147 293 -1127
<< ndcontact >>
rect 517 16 521 26
rect 525 16 529 26
rect 487 5 491 15
rect 495 5 499 15
rect 426 -6 430 4
rect 434 -6 438 4
rect 463 -5 467 5
rect 471 -5 475 5
rect 578 2 582 12
rect 586 2 590 12
rect 487 -20 491 -10
rect 495 -20 499 -10
rect 578 -23 582 -13
rect 586 -23 590 -13
rect -137 -81 -133 -71
rect -129 -81 -125 -71
rect 554 -55 558 -45
rect 562 -55 566 -45
rect -167 -92 -163 -82
rect -159 -92 -155 -82
rect 399 -82 403 -72
rect 407 -82 411 -72
rect -228 -103 -224 -93
rect -220 -103 -216 -93
rect -191 -102 -187 -92
rect -183 -102 -179 -92
rect -76 -95 -72 -85
rect -68 -95 -64 -85
rect -167 -117 -163 -107
rect -159 -117 -155 -107
rect -76 -120 -72 -110
rect -68 -120 -64 -110
rect -100 -152 -96 -142
rect -92 -152 -88 -142
rect -255 -179 -251 -169
rect -247 -179 -243 -169
rect -138 -227 -134 -217
rect -130 -227 -126 -217
rect -168 -238 -164 -228
rect -160 -238 -156 -228
rect -229 -249 -225 -239
rect -221 -249 -217 -239
rect -192 -248 -188 -238
rect -184 -248 -180 -238
rect -77 -241 -73 -231
rect -69 -241 -65 -231
rect -168 -263 -164 -253
rect -160 -263 -156 -253
rect -8 -253 -4 -243
rect 14 -253 18 -243
rect 31 -244 35 -234
rect 53 -244 57 -234
rect -77 -266 -73 -256
rect -69 -266 -65 -256
rect 149 -246 153 -236
rect 171 -246 175 -236
rect 188 -237 192 -227
rect 210 -237 214 -227
rect 517 -244 521 -234
rect 525 -244 529 -234
rect 71 -267 75 -257
rect 93 -267 97 -257
rect 228 -260 232 -250
rect 250 -260 254 -250
rect 487 -255 491 -245
rect 495 -255 499 -245
rect -101 -298 -97 -288
rect -93 -298 -89 -288
rect 426 -266 430 -256
rect 434 -266 438 -256
rect 463 -265 467 -255
rect 471 -265 475 -255
rect 578 -258 582 -248
rect 586 -258 590 -248
rect 31 -313 35 -303
rect 53 -313 57 -303
rect 188 -306 192 -296
rect 210 -306 214 -296
rect 487 -280 491 -270
rect 495 -280 499 -270
rect 578 -283 582 -273
rect 586 -283 590 -273
rect -256 -325 -252 -315
rect -248 -325 -244 -315
rect 554 -315 558 -305
rect 562 -315 566 -305
rect -138 -368 -134 -358
rect -130 -368 -126 -358
rect 399 -342 403 -332
rect 407 -342 411 -332
rect -168 -379 -164 -369
rect -160 -379 -156 -369
rect -229 -390 -225 -380
rect -221 -390 -217 -380
rect -192 -389 -188 -379
rect -184 -389 -180 -379
rect -77 -382 -73 -372
rect -69 -382 -65 -372
rect 24 -379 28 -369
rect 46 -379 50 -369
rect 56 -379 60 -369
rect 68 -379 72 -369
rect -168 -404 -164 -394
rect -160 -404 -156 -394
rect -77 -407 -73 -397
rect -69 -407 -65 -397
rect 140 -403 144 -393
rect 162 -403 166 -393
rect 172 -403 176 -393
rect 184 -403 188 -393
rect 213 -405 217 -395
rect 222 -405 226 -395
rect 231 -405 235 -395
rect 239 -405 243 -395
rect 247 -405 251 -395
rect -101 -439 -97 -429
rect -93 -439 -89 -429
rect -256 -466 -252 -456
rect -248 -466 -244 -456
rect -139 -511 -135 -501
rect -131 -511 -127 -501
rect -169 -522 -165 -512
rect -161 -522 -157 -512
rect -230 -533 -226 -523
rect -222 -533 -218 -523
rect -193 -532 -189 -522
rect -185 -532 -181 -522
rect -78 -525 -74 -515
rect -70 -525 -66 -515
rect -169 -547 -165 -537
rect -161 -547 -157 -537
rect -2 -538 2 -528
rect 20 -538 24 -528
rect 37 -529 41 -519
rect 59 -529 63 -519
rect -78 -550 -74 -540
rect -70 -550 -66 -540
rect 155 -531 159 -521
rect 177 -531 181 -521
rect 194 -522 198 -512
rect 216 -522 220 -512
rect 517 -528 521 -518
rect 525 -528 529 -518
rect 77 -552 81 -542
rect 99 -552 103 -542
rect 234 -545 238 -535
rect 256 -545 260 -535
rect 487 -539 491 -529
rect 495 -539 499 -529
rect -102 -582 -98 -572
rect -94 -582 -90 -572
rect 426 -550 430 -540
rect 434 -550 438 -540
rect 463 -549 467 -539
rect 471 -549 475 -539
rect 578 -542 582 -532
rect 586 -542 590 -532
rect 37 -598 41 -588
rect 59 -598 63 -588
rect 194 -591 198 -581
rect 216 -591 220 -581
rect 487 -564 491 -554
rect 495 -564 499 -554
rect 578 -567 582 -557
rect 586 -567 590 -557
rect -257 -609 -253 -599
rect -249 -609 -245 -599
rect 554 -599 558 -589
rect 562 -599 566 -589
rect -139 -652 -135 -642
rect -131 -652 -127 -642
rect 399 -626 403 -616
rect 407 -626 411 -616
rect -169 -663 -165 -653
rect -161 -663 -157 -653
rect -230 -674 -226 -664
rect -222 -674 -218 -664
rect -193 -673 -189 -663
rect -185 -673 -181 -663
rect -78 -666 -74 -656
rect -70 -666 -66 -656
rect 30 -664 34 -654
rect 52 -664 56 -654
rect 62 -664 66 -654
rect 74 -664 78 -654
rect -169 -688 -165 -678
rect -161 -688 -157 -678
rect -78 -691 -74 -681
rect -70 -691 -66 -681
rect 146 -688 150 -678
rect 168 -688 172 -678
rect 178 -688 182 -678
rect 190 -688 194 -678
rect 219 -688 223 -678
rect 241 -688 245 -678
rect 251 -688 255 -678
rect 263 -688 267 -678
rect 289 -690 293 -680
rect 298 -690 302 -680
rect 307 -690 311 -680
rect 315 -690 319 -680
rect 323 -690 327 -680
rect -102 -723 -98 -713
rect -94 -723 -90 -713
rect -257 -750 -253 -740
rect -249 -750 -245 -740
rect 242 -771 246 -761
rect 251 -771 255 -761
rect 260 -771 264 -761
rect 268 -771 272 -761
rect 276 -771 280 -761
rect -139 -800 -135 -790
rect -131 -800 -127 -790
rect -169 -811 -165 -801
rect -161 -811 -157 -801
rect 517 -797 521 -787
rect 525 -797 529 -787
rect -230 -822 -226 -812
rect -222 -822 -218 -812
rect -193 -821 -189 -811
rect -185 -821 -181 -811
rect -78 -814 -74 -804
rect -70 -814 -66 -804
rect 487 -808 491 -798
rect 495 -808 499 -798
rect -169 -836 -165 -826
rect -161 -836 -157 -826
rect 426 -819 430 -809
rect 434 -819 438 -809
rect 463 -818 467 -808
rect 471 -818 475 -808
rect 578 -811 582 -801
rect 586 -811 590 -801
rect -78 -839 -74 -829
rect -70 -839 -66 -829
rect -102 -871 -98 -861
rect -94 -871 -90 -861
rect 487 -833 491 -823
rect 495 -833 499 -823
rect 578 -836 582 -826
rect 586 -836 590 -826
rect -257 -898 -253 -888
rect -249 -898 -245 -888
rect 554 -868 558 -858
rect 562 -868 566 -858
rect -139 -941 -135 -931
rect -131 -941 -127 -931
rect -2 -918 2 -908
rect 20 -918 24 -908
rect 37 -909 41 -899
rect 59 -909 63 -899
rect 155 -911 159 -901
rect 177 -911 181 -901
rect 194 -902 198 -892
rect 216 -902 220 -892
rect 399 -895 403 -885
rect 407 -895 411 -885
rect 77 -932 81 -922
rect 99 -932 103 -922
rect 234 -925 238 -915
rect 256 -925 260 -915
rect -169 -952 -165 -942
rect -161 -952 -157 -942
rect -230 -963 -226 -953
rect -222 -963 -218 -953
rect -193 -962 -189 -952
rect -185 -962 -181 -952
rect -78 -955 -74 -945
rect -70 -955 -66 -945
rect -169 -977 -165 -967
rect -161 -977 -157 -967
rect -78 -980 -74 -970
rect -70 -980 -66 -970
rect 37 -978 41 -968
rect 59 -978 63 -968
rect 194 -971 198 -961
rect 216 -971 220 -961
rect -102 -1012 -98 -1002
rect -94 -1012 -90 -1002
rect -257 -1039 -253 -1029
rect -249 -1039 -245 -1029
rect 30 -1044 34 -1034
rect 52 -1044 56 -1034
rect 62 -1044 66 -1034
rect 74 -1044 78 -1034
rect 517 -1016 521 -1006
rect 525 -1016 529 -1006
rect 487 -1027 491 -1017
rect 495 -1027 499 -1017
rect 426 -1038 430 -1028
rect 434 -1038 438 -1028
rect 463 -1037 467 -1027
rect 471 -1037 475 -1027
rect 578 -1030 582 -1020
rect 586 -1030 590 -1020
rect 146 -1068 150 -1058
rect 168 -1068 172 -1058
rect 178 -1068 182 -1058
rect 190 -1068 194 -1058
rect 219 -1068 223 -1058
rect 241 -1068 245 -1058
rect 251 -1068 255 -1058
rect 263 -1068 267 -1058
rect 290 -1070 294 -1060
rect 299 -1070 303 -1060
rect 308 -1070 312 -1060
rect 316 -1070 320 -1060
rect 324 -1070 328 -1060
rect 487 -1052 491 -1042
rect 495 -1052 499 -1042
rect 578 -1055 582 -1045
rect 586 -1055 590 -1045
rect 554 -1087 558 -1077
rect 562 -1087 566 -1077
rect 399 -1114 403 -1104
rect 407 -1114 411 -1104
rect 144 -1160 148 -1150
rect 166 -1160 170 -1150
rect 176 -1160 180 -1150
rect 188 -1160 192 -1150
rect 209 -1162 213 -1152
rect 218 -1162 222 -1152
rect 227 -1162 231 -1152
rect 235 -1162 239 -1152
rect 243 -1162 247 -1152
rect 259 -1169 263 -1159
rect 268 -1169 272 -1159
rect 277 -1169 281 -1159
rect 285 -1169 289 -1159
rect 293 -1169 297 -1159
<< pdcontact >>
rect 426 18 430 38
rect 434 18 438 38
rect 487 27 491 47
rect 495 27 499 47
rect 578 24 582 44
rect 586 24 590 44
rect 463 -39 467 -19
rect 471 -39 475 -19
rect 517 -18 521 2
rect 525 -18 529 2
rect 554 -31 558 -11
rect 562 -31 566 -11
rect -228 -79 -224 -59
rect -220 -79 -216 -59
rect -167 -70 -163 -50
rect -159 -70 -155 -50
rect -76 -73 -72 -53
rect -68 -73 -64 -53
rect 399 -60 403 -40
rect 407 -60 411 -40
rect 487 -52 491 -32
rect 495 -52 499 -32
rect 578 -55 582 -35
rect 586 -55 590 -35
rect -191 -136 -187 -116
rect -183 -136 -179 -116
rect -137 -115 -133 -95
rect -129 -115 -125 -95
rect -100 -128 -96 -108
rect -92 -128 -88 -108
rect -255 -157 -251 -137
rect -247 -157 -243 -137
rect -167 -149 -163 -129
rect -159 -149 -155 -129
rect -76 -152 -72 -132
rect -68 -152 -64 -132
rect -229 -225 -225 -205
rect -221 -225 -217 -205
rect -168 -216 -164 -196
rect -160 -216 -156 -196
rect -77 -219 -73 -199
rect -69 -219 -65 -199
rect -8 -228 -4 -208
rect 3 -228 7 -208
rect 14 -228 18 -208
rect 31 -219 35 -199
rect 42 -219 46 -199
rect 53 -219 57 -199
rect -192 -282 -188 -262
rect -184 -282 -180 -262
rect -138 -261 -134 -241
rect -130 -261 -126 -241
rect 149 -221 153 -201
rect 160 -221 164 -201
rect 171 -221 175 -201
rect 188 -212 192 -192
rect 199 -212 203 -192
rect 210 -212 214 -192
rect 71 -242 75 -222
rect 82 -242 86 -222
rect 93 -242 97 -222
rect -101 -274 -97 -254
rect -93 -274 -89 -254
rect 228 -235 232 -215
rect 239 -235 243 -215
rect 250 -235 254 -215
rect 426 -242 430 -222
rect 434 -242 438 -222
rect 487 -233 491 -213
rect 495 -233 499 -213
rect 578 -236 582 -216
rect 586 -236 590 -216
rect -256 -303 -252 -283
rect -248 -303 -244 -283
rect -168 -295 -164 -275
rect -160 -295 -156 -275
rect -77 -298 -73 -278
rect -69 -298 -65 -278
rect 31 -288 35 -268
rect 42 -288 46 -268
rect 53 -288 57 -268
rect 188 -281 192 -261
rect 199 -281 203 -261
rect 210 -281 214 -261
rect 463 -299 467 -279
rect 471 -299 475 -279
rect 517 -278 521 -258
rect 525 -278 529 -258
rect 554 -291 558 -271
rect 562 -291 566 -271
rect 399 -320 403 -300
rect 407 -320 411 -300
rect 487 -312 491 -292
rect 495 -312 499 -292
rect 578 -315 582 -295
rect 586 -315 590 -295
rect -229 -366 -225 -346
rect -221 -366 -217 -346
rect -168 -357 -164 -337
rect -160 -357 -156 -337
rect -77 -360 -73 -340
rect -69 -360 -65 -340
rect 24 -354 28 -334
rect 35 -354 39 -334
rect 46 -354 50 -334
rect 56 -354 60 -334
rect 68 -354 72 -334
rect 140 -378 144 -358
rect 151 -378 155 -358
rect 162 -378 166 -358
rect 172 -378 176 -358
rect 184 -378 188 -358
rect -192 -423 -188 -403
rect -184 -423 -180 -403
rect -138 -402 -134 -382
rect -130 -402 -126 -382
rect 213 -383 217 -363
rect 230 -383 234 -363
rect 239 -383 243 -363
rect 247 -383 251 -363
rect -101 -415 -97 -395
rect -93 -415 -89 -395
rect -256 -444 -252 -424
rect -248 -444 -244 -424
rect -168 -436 -164 -416
rect -160 -436 -156 -416
rect -77 -439 -73 -419
rect -69 -439 -65 -419
rect -230 -509 -226 -489
rect -222 -509 -218 -489
rect -169 -500 -165 -480
rect -161 -500 -157 -480
rect -78 -503 -74 -483
rect -70 -503 -66 -483
rect -2 -513 2 -493
rect 9 -513 13 -493
rect 20 -513 24 -493
rect 37 -504 41 -484
rect 48 -504 52 -484
rect 59 -504 63 -484
rect -193 -566 -189 -546
rect -185 -566 -181 -546
rect -139 -545 -135 -525
rect -131 -545 -127 -525
rect 155 -506 159 -486
rect 166 -506 170 -486
rect 177 -506 181 -486
rect 194 -497 198 -477
rect 205 -497 209 -477
rect 216 -497 220 -477
rect -102 -558 -98 -538
rect -94 -558 -90 -538
rect 77 -527 81 -507
rect 88 -527 92 -507
rect 99 -527 103 -507
rect 234 -520 238 -500
rect 245 -520 249 -500
rect 256 -520 260 -500
rect 426 -526 430 -506
rect 434 -526 438 -506
rect 487 -517 491 -497
rect 495 -517 499 -497
rect 578 -520 582 -500
rect 586 -520 590 -500
rect -257 -587 -253 -567
rect -249 -587 -245 -567
rect -169 -579 -165 -559
rect -161 -579 -157 -559
rect -78 -582 -74 -562
rect -70 -582 -66 -562
rect 37 -573 41 -553
rect 48 -573 52 -553
rect 59 -573 63 -553
rect 194 -566 198 -546
rect 205 -566 209 -546
rect 216 -566 220 -546
rect 463 -583 467 -563
rect 471 -583 475 -563
rect 517 -562 521 -542
rect 525 -562 529 -542
rect 554 -575 558 -555
rect 562 -575 566 -555
rect 399 -604 403 -584
rect 407 -604 411 -584
rect 487 -596 491 -576
rect 495 -596 499 -576
rect 578 -599 582 -579
rect 586 -599 590 -579
rect -230 -650 -226 -630
rect -222 -650 -218 -630
rect -169 -641 -165 -621
rect -161 -641 -157 -621
rect -78 -644 -74 -624
rect -70 -644 -66 -624
rect 30 -639 34 -619
rect 41 -639 45 -619
rect 52 -639 56 -619
rect 62 -639 66 -619
rect 74 -639 78 -619
rect 146 -663 150 -643
rect 157 -663 161 -643
rect 168 -663 172 -643
rect 178 -663 182 -643
rect 190 -663 194 -643
rect 219 -663 223 -643
rect 230 -663 234 -643
rect 241 -663 245 -643
rect 251 -663 255 -643
rect 263 -663 267 -643
rect -193 -707 -189 -687
rect -185 -707 -181 -687
rect -139 -686 -135 -666
rect -131 -686 -127 -666
rect 289 -668 293 -648
rect 306 -668 310 -648
rect 315 -668 319 -648
rect 323 -668 327 -648
rect -102 -699 -98 -679
rect -94 -699 -90 -679
rect -257 -728 -253 -708
rect -249 -728 -245 -708
rect -169 -720 -165 -700
rect -161 -720 -157 -700
rect -78 -723 -74 -703
rect -70 -723 -66 -703
rect 242 -749 246 -729
rect 259 -749 263 -729
rect 268 -749 272 -729
rect 276 -749 280 -729
rect -230 -798 -226 -778
rect -222 -798 -218 -778
rect -169 -789 -165 -769
rect -161 -789 -157 -769
rect -78 -792 -74 -772
rect -70 -792 -66 -772
rect 426 -795 430 -775
rect 434 -795 438 -775
rect 487 -786 491 -766
rect 495 -786 499 -766
rect 578 -789 582 -769
rect 586 -789 590 -769
rect -193 -855 -189 -835
rect -185 -855 -181 -835
rect -139 -834 -135 -814
rect -131 -834 -127 -814
rect -102 -847 -98 -827
rect -94 -847 -90 -827
rect -257 -876 -253 -856
rect -249 -876 -245 -856
rect -169 -868 -165 -848
rect -161 -868 -157 -848
rect -78 -871 -74 -851
rect -70 -871 -66 -851
rect 463 -852 467 -832
rect 471 -852 475 -832
rect 517 -831 521 -811
rect 525 -831 529 -811
rect 554 -844 558 -824
rect 562 -844 566 -824
rect -2 -893 2 -873
rect 9 -893 13 -873
rect 20 -893 24 -873
rect 37 -884 41 -864
rect 48 -884 52 -864
rect 59 -884 63 -864
rect 155 -886 159 -866
rect 166 -886 170 -866
rect 177 -886 181 -866
rect 194 -877 198 -857
rect 205 -877 209 -857
rect 216 -877 220 -857
rect 399 -873 403 -853
rect 407 -873 411 -853
rect 487 -865 491 -845
rect 495 -865 499 -845
rect 578 -868 582 -848
rect 586 -868 590 -848
rect -230 -939 -226 -919
rect -222 -939 -218 -919
rect -169 -930 -165 -910
rect -161 -930 -157 -910
rect -78 -933 -74 -913
rect -70 -933 -66 -913
rect 77 -907 81 -887
rect 88 -907 92 -887
rect 99 -907 103 -887
rect 234 -900 238 -880
rect 245 -900 249 -880
rect 256 -900 260 -880
rect 37 -953 41 -933
rect 48 -953 52 -933
rect 59 -953 63 -933
rect 194 -946 198 -926
rect 205 -946 209 -926
rect 216 -946 220 -926
rect -193 -996 -189 -976
rect -185 -996 -181 -976
rect -139 -975 -135 -955
rect -131 -975 -127 -955
rect -102 -988 -98 -968
rect -94 -988 -90 -968
rect -257 -1017 -253 -997
rect -249 -1017 -245 -997
rect -169 -1009 -165 -989
rect -161 -1009 -157 -989
rect -78 -1012 -74 -992
rect -70 -1012 -66 -992
rect 30 -1019 34 -999
rect 41 -1019 45 -999
rect 52 -1019 56 -999
rect 62 -1019 66 -999
rect 74 -1019 78 -999
rect 426 -1014 430 -994
rect 434 -1014 438 -994
rect 487 -1005 491 -985
rect 495 -1005 499 -985
rect 146 -1043 150 -1023
rect 157 -1043 161 -1023
rect 168 -1043 172 -1023
rect 178 -1043 182 -1023
rect 190 -1043 194 -1023
rect 219 -1043 223 -1023
rect 230 -1043 234 -1023
rect 241 -1043 245 -1023
rect 251 -1043 255 -1023
rect 263 -1043 267 -1023
rect 578 -1008 582 -988
rect 586 -1008 590 -988
rect 290 -1048 294 -1028
rect 307 -1048 311 -1028
rect 316 -1048 320 -1028
rect 324 -1048 328 -1028
rect 463 -1071 467 -1051
rect 471 -1071 475 -1051
rect 517 -1050 521 -1030
rect 525 -1050 529 -1030
rect 554 -1063 558 -1043
rect 562 -1063 566 -1043
rect 399 -1092 403 -1072
rect 407 -1092 411 -1072
rect 487 -1084 491 -1064
rect 495 -1084 499 -1064
rect 578 -1087 582 -1067
rect 586 -1087 590 -1067
rect 144 -1135 148 -1115
rect 155 -1135 159 -1115
rect 166 -1135 170 -1115
rect 176 -1135 180 -1115
rect 188 -1135 192 -1115
rect 209 -1140 213 -1120
rect 226 -1140 230 -1120
rect 235 -1140 239 -1120
rect 243 -1140 247 -1120
rect 259 -1147 263 -1127
rect 276 -1147 280 -1127
rect 285 -1147 289 -1127
rect 293 -1147 297 -1127
<< polysilicon >>
rect 492 47 494 50
rect 431 38 433 45
rect 583 44 585 47
rect 431 13 433 18
rect 492 15 494 27
rect 522 26 524 33
rect 431 4 433 9
rect 468 5 470 12
rect 522 11 524 16
rect 583 12 585 24
rect 492 2 494 5
rect 522 2 524 7
rect 431 -13 433 -6
rect 468 -10 470 -5
rect 492 -10 494 -7
rect 468 -19 470 -14
rect 404 -40 406 -37
rect 583 -1 585 2
rect 559 -11 561 -4
rect 492 -32 494 -20
rect 522 -25 524 -18
rect 583 -13 585 -10
rect -162 -50 -160 -47
rect -223 -59 -221 -52
rect -71 -53 -69 -50
rect -223 -84 -221 -79
rect -162 -82 -160 -70
rect -132 -71 -130 -64
rect 468 -46 470 -39
rect 559 -36 561 -31
rect 583 -35 585 -23
rect 559 -45 561 -40
rect 492 -55 494 -52
rect 404 -72 406 -60
rect 559 -62 561 -55
rect 583 -58 585 -55
rect -223 -93 -221 -88
rect -186 -92 -184 -85
rect -132 -86 -130 -81
rect -71 -85 -69 -73
rect 98 -77 100 -76
rect 105 -77 107 -76
rect 404 -85 406 -82
rect -162 -95 -160 -92
rect -132 -95 -130 -90
rect -223 -110 -221 -103
rect -186 -107 -184 -102
rect -162 -107 -160 -104
rect -186 -116 -184 -111
rect -250 -137 -248 -134
rect -71 -98 -69 -95
rect -95 -108 -93 -101
rect -162 -129 -160 -117
rect -132 -122 -130 -115
rect -71 -110 -69 -107
rect -186 -143 -184 -136
rect -95 -133 -93 -128
rect -71 -132 -69 -120
rect -95 -142 -93 -137
rect -162 -152 -160 -149
rect -250 -169 -248 -157
rect -95 -159 -93 -152
rect -71 -155 -69 -152
rect -250 -182 -248 -179
rect 193 -192 195 -189
rect 207 -192 209 -189
rect -163 -196 -161 -193
rect -224 -205 -222 -198
rect -72 -199 -70 -196
rect 36 -199 38 -196
rect 50 -199 52 -196
rect -224 -230 -222 -225
rect -163 -228 -161 -216
rect -133 -217 -131 -210
rect -3 -208 -1 -205
rect 11 -208 13 -205
rect -224 -239 -222 -234
rect -187 -238 -185 -231
rect -133 -232 -131 -227
rect -72 -231 -70 -219
rect 154 -201 156 -198
rect 168 -201 170 -198
rect -163 -241 -161 -238
rect -133 -241 -131 -236
rect -224 -256 -222 -249
rect -187 -253 -185 -248
rect -163 -253 -161 -250
rect -187 -262 -185 -257
rect -251 -283 -249 -280
rect -72 -244 -70 -241
rect -3 -243 -1 -228
rect 11 -243 13 -228
rect 36 -234 38 -219
rect 50 -234 52 -219
rect 76 -222 78 -219
rect 90 -222 92 -219
rect -96 -254 -94 -247
rect 154 -236 156 -221
rect 168 -236 170 -221
rect 193 -227 195 -212
rect 207 -227 209 -212
rect 233 -215 235 -212
rect 247 -215 249 -212
rect 492 -213 494 -210
rect 36 -249 38 -244
rect 50 -249 52 -244
rect -163 -275 -161 -263
rect -133 -268 -131 -261
rect -72 -256 -70 -253
rect -3 -258 -1 -253
rect 11 -258 13 -253
rect 76 -257 78 -242
rect 90 -257 92 -242
rect 431 -222 433 -215
rect 193 -242 195 -237
rect 207 -242 209 -237
rect 154 -251 156 -246
rect 168 -251 170 -246
rect 233 -250 235 -235
rect 247 -250 249 -235
rect 583 -216 585 -213
rect 431 -247 433 -242
rect 492 -245 494 -233
rect 522 -234 524 -227
rect -187 -289 -185 -282
rect -96 -279 -94 -274
rect -72 -278 -70 -266
rect 36 -268 38 -265
rect 50 -268 52 -265
rect 193 -261 195 -258
rect 207 -261 209 -258
rect 431 -256 433 -251
rect 468 -255 470 -248
rect 522 -249 524 -244
rect 583 -248 585 -236
rect -96 -288 -94 -283
rect -163 -298 -161 -295
rect 76 -272 78 -267
rect 90 -272 92 -267
rect 233 -265 235 -260
rect 247 -265 249 -260
rect 492 -258 494 -255
rect 522 -258 524 -253
rect 431 -273 433 -266
rect 468 -270 470 -265
rect 492 -270 494 -267
rect 468 -279 470 -274
rect -251 -315 -249 -303
rect -96 -305 -94 -298
rect -72 -301 -70 -298
rect 36 -303 38 -288
rect 50 -303 52 -288
rect 193 -296 195 -281
rect 207 -296 209 -281
rect 404 -300 406 -297
rect 583 -261 585 -258
rect 559 -271 561 -264
rect 492 -292 494 -280
rect 522 -285 524 -278
rect 583 -273 585 -270
rect 193 -311 195 -306
rect 207 -311 209 -306
rect 36 -318 38 -313
rect 50 -318 52 -313
rect 468 -306 470 -299
rect 559 -296 561 -291
rect 583 -295 585 -283
rect 559 -305 561 -300
rect 492 -315 494 -312
rect -251 -328 -249 -325
rect 29 -334 31 -331
rect 43 -334 45 -331
rect 63 -334 65 -331
rect 404 -332 406 -320
rect 559 -322 561 -315
rect 583 -318 585 -315
rect -163 -337 -161 -334
rect -224 -346 -222 -339
rect -72 -340 -70 -337
rect -224 -371 -222 -366
rect -163 -369 -161 -357
rect -133 -358 -131 -351
rect 404 -345 406 -342
rect -224 -380 -222 -375
rect -187 -379 -185 -372
rect -133 -373 -131 -368
rect -72 -372 -70 -360
rect 29 -369 31 -354
rect 43 -369 45 -354
rect 63 -369 65 -354
rect 145 -358 147 -355
rect 159 -358 161 -355
rect 179 -358 181 -355
rect -163 -382 -161 -379
rect -133 -382 -131 -377
rect 219 -363 221 -349
rect 226 -363 228 -349
rect 244 -363 246 -360
rect -224 -397 -222 -390
rect -187 -394 -185 -389
rect -163 -394 -161 -391
rect -187 -403 -185 -398
rect -251 -424 -249 -421
rect -72 -385 -70 -382
rect 29 -384 31 -379
rect 43 -384 45 -379
rect 63 -382 65 -379
rect -96 -395 -94 -388
rect 145 -393 147 -378
rect 159 -393 161 -378
rect 179 -393 181 -378
rect -163 -416 -161 -404
rect -133 -409 -131 -402
rect -72 -397 -70 -394
rect 219 -395 221 -383
rect 226 -391 228 -383
rect 226 -393 229 -391
rect 227 -395 229 -393
rect 244 -395 246 -383
rect -187 -430 -185 -423
rect -96 -420 -94 -415
rect -72 -419 -70 -407
rect 145 -408 147 -403
rect 159 -408 161 -403
rect 179 -406 181 -403
rect 219 -408 221 -405
rect 227 -408 229 -405
rect 244 -408 246 -405
rect -96 -429 -94 -424
rect -163 -439 -161 -436
rect -251 -456 -249 -444
rect -96 -446 -94 -439
rect -72 -442 -70 -439
rect -251 -469 -249 -466
rect 199 -477 201 -474
rect 213 -477 215 -474
rect -164 -480 -162 -477
rect -225 -489 -223 -482
rect -73 -483 -71 -480
rect -225 -514 -223 -509
rect -164 -512 -162 -500
rect -134 -501 -132 -494
rect 42 -484 44 -481
rect 56 -484 58 -481
rect 3 -493 5 -490
rect 17 -493 19 -490
rect -225 -523 -223 -518
rect -188 -522 -186 -515
rect -134 -516 -132 -511
rect -73 -515 -71 -503
rect 160 -486 162 -483
rect 174 -486 176 -483
rect -164 -525 -162 -522
rect -134 -525 -132 -520
rect -225 -540 -223 -533
rect -188 -537 -186 -532
rect -164 -537 -162 -534
rect -188 -546 -186 -541
rect -252 -567 -250 -564
rect -73 -528 -71 -525
rect 3 -528 5 -513
rect 17 -528 19 -513
rect 42 -519 44 -504
rect 56 -519 58 -504
rect 82 -507 84 -504
rect 96 -507 98 -504
rect 492 -497 494 -494
rect -97 -538 -95 -531
rect -164 -559 -162 -547
rect -134 -552 -132 -545
rect -73 -540 -71 -537
rect 160 -521 162 -506
rect 174 -521 176 -506
rect 199 -512 201 -497
rect 213 -512 215 -497
rect 239 -500 241 -497
rect 253 -500 255 -497
rect 42 -534 44 -529
rect 56 -534 58 -529
rect 3 -543 5 -538
rect 17 -543 19 -538
rect 82 -542 84 -527
rect 96 -542 98 -527
rect 431 -506 433 -499
rect 199 -527 201 -522
rect 213 -527 215 -522
rect 160 -536 162 -531
rect 174 -536 176 -531
rect 239 -535 241 -520
rect 253 -535 255 -520
rect 583 -500 585 -497
rect 431 -531 433 -526
rect 492 -529 494 -517
rect 522 -518 524 -511
rect -188 -573 -186 -566
rect -97 -563 -95 -558
rect -73 -562 -71 -550
rect 42 -553 44 -550
rect 56 -553 58 -550
rect 199 -546 201 -543
rect 213 -546 215 -543
rect 431 -540 433 -535
rect 468 -539 470 -532
rect 522 -533 524 -528
rect 583 -532 585 -520
rect -97 -572 -95 -567
rect -164 -582 -162 -579
rect 82 -557 84 -552
rect 96 -557 98 -552
rect 239 -550 241 -545
rect 253 -550 255 -545
rect 492 -542 494 -539
rect 522 -542 524 -537
rect 431 -557 433 -550
rect 468 -554 470 -549
rect 492 -554 494 -551
rect 468 -563 470 -558
rect -252 -599 -250 -587
rect -97 -589 -95 -582
rect -73 -585 -71 -582
rect 42 -588 44 -573
rect 56 -588 58 -573
rect 199 -581 201 -566
rect 213 -581 215 -566
rect 404 -584 406 -581
rect 583 -545 585 -542
rect 559 -555 561 -548
rect 492 -576 494 -564
rect 522 -569 524 -562
rect 583 -557 585 -554
rect 199 -596 201 -591
rect 213 -596 215 -591
rect 42 -603 44 -598
rect 56 -603 58 -598
rect 468 -590 470 -583
rect 559 -580 561 -575
rect 583 -579 585 -567
rect 559 -589 561 -584
rect 492 -599 494 -596
rect -252 -612 -250 -609
rect 404 -616 406 -604
rect 559 -606 561 -599
rect 583 -602 585 -599
rect -164 -621 -162 -618
rect 35 -619 37 -616
rect 49 -619 51 -616
rect 69 -619 71 -616
rect -225 -630 -223 -623
rect -73 -624 -71 -621
rect -225 -655 -223 -650
rect -164 -653 -162 -641
rect -134 -642 -132 -635
rect 404 -629 406 -626
rect -225 -664 -223 -659
rect -188 -663 -186 -656
rect -134 -657 -132 -652
rect -73 -656 -71 -644
rect 35 -654 37 -639
rect 49 -654 51 -639
rect 69 -654 71 -639
rect 151 -643 153 -640
rect 165 -643 167 -640
rect 185 -643 187 -640
rect 224 -643 226 -640
rect 238 -643 240 -640
rect 258 -643 260 -640
rect -164 -666 -162 -663
rect -134 -666 -132 -661
rect 295 -648 297 -634
rect 302 -648 304 -634
rect 320 -648 322 -645
rect -225 -681 -223 -674
rect -188 -678 -186 -673
rect -164 -678 -162 -675
rect -188 -687 -186 -682
rect -252 -708 -250 -705
rect -73 -669 -71 -666
rect 35 -669 37 -664
rect 49 -669 51 -664
rect 69 -667 71 -664
rect -97 -679 -95 -672
rect 151 -678 153 -663
rect 165 -678 167 -663
rect 185 -678 187 -663
rect 224 -678 226 -663
rect 238 -678 240 -663
rect 258 -678 260 -663
rect -164 -700 -162 -688
rect -134 -693 -132 -686
rect -73 -681 -71 -678
rect 295 -680 297 -668
rect 302 -676 304 -668
rect 302 -678 305 -676
rect 303 -680 305 -678
rect 320 -680 322 -668
rect -188 -714 -186 -707
rect -97 -704 -95 -699
rect -73 -703 -71 -691
rect 151 -693 153 -688
rect 165 -693 167 -688
rect 185 -691 187 -688
rect 224 -693 226 -688
rect 238 -693 240 -688
rect 258 -691 260 -688
rect 295 -693 297 -690
rect 303 -693 305 -690
rect 320 -693 322 -690
rect -97 -713 -95 -708
rect -164 -723 -162 -720
rect -252 -740 -250 -728
rect -97 -730 -95 -723
rect -73 -726 -71 -723
rect 248 -729 250 -715
rect 255 -729 257 -715
rect 273 -729 275 -726
rect -252 -753 -250 -750
rect 248 -761 250 -749
rect 255 -757 257 -749
rect 255 -759 258 -757
rect 256 -761 258 -759
rect 273 -761 275 -749
rect -164 -769 -162 -766
rect -225 -778 -223 -771
rect -73 -772 -71 -769
rect 492 -766 494 -763
rect -225 -803 -223 -798
rect -164 -801 -162 -789
rect -134 -790 -132 -783
rect 248 -774 250 -771
rect 256 -774 258 -771
rect 273 -774 275 -771
rect 431 -775 433 -768
rect -225 -812 -223 -807
rect -188 -811 -186 -804
rect -134 -805 -132 -800
rect -73 -804 -71 -792
rect 583 -769 585 -766
rect 431 -800 433 -795
rect 492 -798 494 -786
rect 522 -787 524 -780
rect -164 -814 -162 -811
rect -134 -814 -132 -809
rect 431 -809 433 -804
rect 468 -808 470 -801
rect 522 -802 524 -797
rect 583 -801 585 -789
rect -225 -829 -223 -822
rect -188 -826 -186 -821
rect -164 -826 -162 -823
rect -188 -835 -186 -830
rect -252 -856 -250 -853
rect -73 -817 -71 -814
rect 492 -811 494 -808
rect 522 -811 524 -806
rect -97 -827 -95 -820
rect 431 -826 433 -819
rect 468 -823 470 -818
rect 492 -823 494 -820
rect -164 -848 -162 -836
rect -134 -841 -132 -834
rect -73 -829 -71 -826
rect 468 -832 470 -827
rect -188 -862 -186 -855
rect -97 -852 -95 -847
rect -73 -851 -71 -839
rect -97 -861 -95 -856
rect -164 -871 -162 -868
rect 404 -853 406 -850
rect 583 -814 585 -811
rect 559 -824 561 -817
rect 492 -845 494 -833
rect 522 -838 524 -831
rect 583 -826 585 -823
rect 199 -857 201 -854
rect 213 -857 215 -854
rect 42 -864 44 -861
rect 56 -864 58 -861
rect -252 -888 -250 -876
rect -97 -878 -95 -871
rect -73 -874 -71 -871
rect 3 -873 5 -870
rect 17 -873 19 -870
rect 160 -866 162 -863
rect 174 -866 176 -863
rect -252 -901 -250 -898
rect -164 -910 -162 -907
rect 3 -908 5 -893
rect 17 -908 19 -893
rect 42 -899 44 -884
rect 56 -899 58 -884
rect 82 -887 84 -884
rect 96 -887 98 -884
rect 468 -859 470 -852
rect 559 -849 561 -844
rect 583 -848 585 -836
rect 559 -858 561 -853
rect 492 -868 494 -865
rect -225 -919 -223 -912
rect -73 -913 -71 -910
rect -225 -944 -223 -939
rect -164 -942 -162 -930
rect -134 -931 -132 -924
rect 160 -901 162 -886
rect 174 -901 176 -886
rect 199 -892 201 -877
rect 213 -892 215 -877
rect 239 -880 241 -877
rect 253 -880 255 -877
rect 42 -914 44 -909
rect 56 -914 58 -909
rect 3 -923 5 -918
rect 17 -923 19 -918
rect 82 -922 84 -907
rect 96 -922 98 -907
rect 404 -885 406 -873
rect 559 -875 561 -868
rect 583 -871 585 -868
rect 404 -898 406 -895
rect 199 -906 201 -902
rect 213 -907 215 -902
rect 160 -916 162 -911
rect 174 -916 176 -911
rect 239 -915 241 -900
rect 253 -915 255 -900
rect 42 -933 44 -930
rect 56 -933 58 -930
rect 199 -926 201 -923
rect 213 -926 215 -923
rect -225 -953 -223 -948
rect -188 -952 -186 -945
rect -134 -946 -132 -941
rect -73 -945 -71 -933
rect -164 -955 -162 -952
rect -134 -955 -132 -950
rect 82 -937 84 -932
rect 96 -937 98 -932
rect 239 -930 241 -925
rect 253 -930 255 -925
rect -225 -970 -223 -963
rect -188 -967 -186 -962
rect -164 -967 -162 -964
rect -188 -976 -186 -971
rect -252 -997 -250 -994
rect -73 -958 -71 -955
rect -97 -968 -95 -961
rect -164 -989 -162 -977
rect -134 -982 -132 -975
rect -73 -970 -71 -967
rect 42 -968 44 -953
rect 56 -968 58 -953
rect 199 -961 201 -946
rect 213 -961 215 -946
rect 199 -976 201 -971
rect 213 -976 215 -971
rect -188 -1003 -186 -996
rect -97 -993 -95 -988
rect -73 -992 -71 -980
rect 42 -983 44 -978
rect 56 -983 58 -978
rect 492 -985 494 -982
rect -97 -1002 -95 -997
rect -164 -1012 -162 -1009
rect 431 -994 433 -987
rect 35 -999 37 -996
rect 49 -999 51 -996
rect 69 -999 71 -996
rect -252 -1029 -250 -1017
rect -97 -1019 -95 -1012
rect -73 -1015 -71 -1012
rect 583 -988 585 -985
rect 35 -1034 37 -1019
rect 49 -1034 51 -1019
rect 69 -1034 71 -1019
rect 151 -1023 153 -1020
rect 165 -1023 167 -1020
rect 185 -1023 187 -1020
rect 224 -1023 226 -1020
rect 238 -1023 240 -1020
rect 258 -1023 260 -1020
rect -252 -1042 -250 -1039
rect 296 -1028 298 -1014
rect 303 -1028 305 -1014
rect 431 -1019 433 -1014
rect 492 -1017 494 -1005
rect 522 -1006 524 -999
rect 321 -1028 323 -1025
rect 431 -1028 433 -1023
rect 468 -1027 470 -1020
rect 522 -1021 524 -1016
rect 583 -1020 585 -1008
rect 35 -1049 37 -1044
rect 49 -1049 51 -1044
rect 69 -1047 71 -1044
rect 151 -1058 153 -1043
rect 165 -1058 167 -1043
rect 185 -1058 187 -1043
rect 224 -1058 226 -1043
rect 238 -1058 240 -1043
rect 258 -1058 260 -1043
rect 492 -1030 494 -1027
rect 522 -1030 524 -1025
rect 431 -1045 433 -1038
rect 468 -1042 470 -1037
rect 492 -1042 494 -1039
rect 296 -1060 298 -1048
rect 303 -1056 305 -1048
rect 303 -1058 306 -1056
rect 304 -1060 306 -1058
rect 321 -1060 323 -1048
rect 468 -1051 470 -1046
rect 151 -1073 153 -1068
rect 165 -1073 167 -1068
rect 185 -1071 187 -1068
rect 224 -1073 226 -1068
rect 238 -1073 240 -1068
rect 258 -1071 260 -1068
rect 296 -1073 298 -1070
rect 304 -1073 306 -1070
rect 321 -1073 323 -1070
rect 404 -1072 406 -1069
rect 583 -1033 585 -1030
rect 559 -1043 561 -1036
rect 492 -1064 494 -1052
rect 522 -1057 524 -1050
rect 583 -1045 585 -1042
rect 468 -1078 470 -1071
rect 559 -1068 561 -1063
rect 583 -1067 585 -1055
rect 559 -1077 561 -1072
rect 492 -1087 494 -1084
rect 404 -1104 406 -1092
rect 559 -1094 561 -1087
rect 583 -1090 585 -1087
rect 149 -1115 151 -1112
rect 163 -1115 165 -1112
rect 183 -1115 185 -1112
rect 215 -1120 217 -1106
rect 222 -1120 224 -1106
rect 240 -1120 242 -1117
rect 149 -1150 151 -1135
rect 163 -1150 165 -1135
rect 183 -1150 185 -1135
rect 265 -1127 267 -1113
rect 272 -1127 274 -1113
rect 404 -1117 406 -1114
rect 290 -1127 292 -1124
rect 215 -1152 217 -1140
rect 222 -1148 224 -1140
rect 222 -1150 225 -1148
rect 223 -1152 225 -1150
rect 240 -1152 242 -1140
rect 149 -1165 151 -1160
rect 163 -1165 165 -1160
rect 183 -1163 185 -1160
rect 265 -1159 267 -1147
rect 272 -1155 274 -1147
rect 272 -1157 275 -1155
rect 273 -1159 275 -1157
rect 290 -1159 292 -1147
rect 215 -1165 217 -1162
rect 223 -1165 225 -1162
rect 240 -1165 242 -1162
rect 265 -1172 267 -1169
rect 273 -1172 275 -1169
rect 290 -1172 292 -1169
<< polycontact >>
rect 427 41 431 45
rect 518 29 522 33
rect 488 20 492 24
rect 579 17 583 21
rect 464 8 468 12
rect 427 -13 431 -9
rect 555 -8 559 -4
rect 518 -25 522 -21
rect 494 -29 498 -25
rect -227 -56 -223 -52
rect -136 -68 -132 -64
rect -166 -77 -162 -73
rect 464 -46 468 -42
rect 585 -32 589 -28
rect 400 -67 404 -63
rect 555 -62 559 -58
rect -75 -80 -71 -76
rect -190 -89 -186 -85
rect 94 -80 98 -76
rect 107 -80 111 -76
rect -227 -110 -223 -106
rect -99 -105 -95 -101
rect -136 -122 -132 -118
rect -160 -126 -156 -122
rect -190 -143 -186 -139
rect -69 -129 -65 -125
rect -254 -164 -250 -160
rect -99 -159 -95 -155
rect -228 -202 -224 -198
rect -137 -214 -133 -210
rect -167 -223 -163 -219
rect -76 -226 -72 -222
rect -191 -235 -187 -231
rect -228 -256 -224 -252
rect 32 -230 36 -226
rect -100 -251 -96 -247
rect 189 -223 193 -219
rect 46 -249 50 -245
rect 72 -251 76 -247
rect -137 -268 -133 -264
rect -161 -272 -157 -268
rect -1 -258 3 -254
rect 7 -258 11 -254
rect 86 -256 90 -252
rect 427 -219 431 -215
rect 203 -242 207 -238
rect 229 -244 233 -240
rect 156 -251 160 -247
rect 164 -251 168 -247
rect 243 -249 247 -245
rect 518 -231 522 -227
rect 488 -240 492 -236
rect 579 -243 583 -239
rect -191 -289 -187 -285
rect 464 -252 468 -248
rect -70 -275 -66 -271
rect 427 -273 431 -269
rect 32 -297 36 -293
rect -255 -310 -251 -306
rect -100 -305 -96 -301
rect 189 -290 193 -286
rect 555 -268 559 -264
rect 518 -285 522 -281
rect 494 -289 498 -285
rect 203 -311 207 -307
rect 46 -318 50 -314
rect 464 -306 468 -302
rect 585 -292 589 -288
rect 400 -327 404 -323
rect 555 -322 559 -318
rect -228 -343 -224 -339
rect -137 -355 -133 -351
rect -167 -364 -163 -360
rect 215 -353 219 -349
rect -76 -367 -72 -363
rect -191 -376 -187 -372
rect 25 -366 29 -362
rect 39 -368 43 -364
rect 59 -361 63 -357
rect 228 -353 232 -349
rect -228 -397 -224 -393
rect -100 -392 -96 -388
rect 141 -390 145 -386
rect 155 -392 159 -388
rect 175 -385 179 -381
rect -137 -409 -133 -405
rect -161 -413 -157 -409
rect 240 -390 244 -386
rect -191 -430 -187 -426
rect -70 -416 -66 -412
rect -255 -451 -251 -447
rect -100 -446 -96 -442
rect -229 -486 -225 -482
rect -138 -498 -134 -494
rect -168 -507 -164 -503
rect -77 -510 -73 -506
rect -192 -519 -188 -515
rect -229 -540 -225 -536
rect 38 -515 42 -511
rect -101 -535 -97 -531
rect -138 -552 -134 -548
rect -162 -556 -158 -552
rect 195 -508 199 -504
rect 52 -534 56 -530
rect 78 -536 82 -532
rect 5 -543 9 -539
rect 13 -543 17 -539
rect 92 -541 96 -537
rect 427 -503 431 -499
rect 209 -527 213 -523
rect 235 -529 239 -525
rect 162 -536 166 -532
rect 170 -536 174 -532
rect 249 -534 253 -530
rect 518 -515 522 -511
rect 488 -524 492 -520
rect 579 -527 583 -523
rect -192 -573 -188 -569
rect 464 -536 468 -532
rect -71 -559 -67 -555
rect 427 -557 431 -553
rect 38 -582 42 -578
rect -256 -594 -252 -590
rect -101 -589 -97 -585
rect 195 -575 199 -571
rect 555 -552 559 -548
rect 518 -569 522 -565
rect 494 -573 498 -569
rect 209 -596 213 -592
rect 52 -603 56 -599
rect 464 -590 468 -586
rect 585 -576 589 -572
rect 400 -611 404 -607
rect 555 -606 559 -602
rect -229 -627 -225 -623
rect -138 -639 -134 -635
rect -168 -648 -164 -644
rect 291 -638 295 -634
rect -77 -651 -73 -647
rect -192 -660 -188 -656
rect 31 -651 35 -647
rect 45 -653 49 -649
rect 65 -646 69 -642
rect 304 -638 308 -634
rect -229 -681 -225 -677
rect -101 -676 -97 -672
rect 147 -675 151 -671
rect 161 -677 165 -673
rect 181 -670 185 -666
rect 220 -675 224 -671
rect 234 -677 238 -673
rect 254 -670 258 -666
rect -138 -693 -134 -689
rect -162 -697 -158 -693
rect 316 -675 320 -671
rect -192 -714 -188 -710
rect -71 -700 -67 -696
rect 244 -719 248 -715
rect -256 -735 -252 -731
rect -101 -730 -97 -726
rect 257 -719 261 -715
rect 269 -756 273 -752
rect -229 -775 -225 -771
rect -138 -787 -134 -783
rect -168 -796 -164 -792
rect 427 -772 431 -768
rect -77 -799 -73 -795
rect -192 -808 -188 -804
rect 518 -784 522 -780
rect 488 -793 492 -789
rect 579 -796 583 -792
rect 464 -805 468 -801
rect -229 -829 -225 -825
rect -101 -824 -97 -820
rect 427 -826 431 -822
rect -138 -841 -134 -837
rect -162 -845 -158 -841
rect -192 -862 -188 -858
rect -71 -848 -67 -844
rect 555 -821 559 -817
rect 518 -838 522 -834
rect 494 -842 498 -838
rect -256 -883 -252 -879
rect -101 -878 -97 -874
rect 38 -895 42 -891
rect 464 -859 468 -855
rect 585 -845 589 -841
rect -229 -916 -225 -912
rect -138 -928 -134 -924
rect -168 -937 -164 -933
rect 195 -888 199 -884
rect 400 -880 404 -876
rect 52 -914 56 -910
rect 78 -916 82 -912
rect 5 -923 9 -919
rect 13 -923 17 -919
rect 92 -921 96 -917
rect 555 -875 559 -871
rect 209 -907 213 -903
rect 235 -909 239 -905
rect 162 -916 166 -912
rect 170 -916 174 -912
rect 249 -914 253 -910
rect -77 -940 -73 -936
rect -192 -949 -188 -945
rect -229 -970 -225 -966
rect -101 -965 -97 -961
rect 38 -962 42 -958
rect -138 -982 -134 -978
rect -162 -986 -158 -982
rect 195 -955 199 -951
rect 209 -976 213 -972
rect -192 -1003 -188 -999
rect 52 -983 56 -979
rect -71 -989 -67 -985
rect 427 -991 431 -987
rect -256 -1024 -252 -1020
rect -101 -1019 -97 -1015
rect 518 -1003 522 -999
rect 488 -1012 492 -1008
rect 292 -1018 296 -1014
rect 31 -1031 35 -1027
rect 45 -1033 49 -1029
rect 65 -1026 69 -1022
rect 305 -1018 309 -1014
rect 579 -1015 583 -1011
rect 464 -1024 468 -1020
rect 147 -1055 151 -1051
rect 161 -1057 165 -1053
rect 181 -1050 185 -1046
rect 220 -1055 224 -1051
rect 234 -1057 238 -1053
rect 254 -1050 258 -1046
rect 427 -1045 431 -1041
rect 317 -1055 321 -1051
rect 555 -1040 559 -1036
rect 518 -1057 522 -1053
rect 494 -1061 498 -1057
rect 464 -1078 468 -1074
rect 585 -1064 589 -1060
rect 400 -1099 404 -1095
rect 555 -1094 559 -1090
rect 211 -1110 215 -1106
rect 224 -1110 228 -1106
rect 261 -1117 265 -1113
rect 145 -1147 149 -1143
rect 159 -1149 163 -1145
rect 179 -1142 183 -1138
rect 274 -1117 278 -1113
rect 236 -1147 240 -1143
rect 286 -1154 290 -1150
<< metal1 >>
rect -278 88 -275 100
rect -170 99 -162 101
rect -79 96 -71 98
rect -278 85 -229 88
rect -296 62 -292 65
rect -278 57 -275 85
rect 229 65 234 67
rect -242 57 -239 61
rect 39 58 43 62
rect -53 52 -49 55
rect -278 -19 -275 52
rect -169 40 -167 43
rect -78 37 -75 40
rect -52 37 -49 52
rect 103 50 174 53
rect -52 34 -20 37
rect -47 25 -29 28
rect -258 12 -250 14
rect -152 -16 -150 -13
rect -61 -19 -59 -16
rect -278 -23 -260 -19
rect -278 -53 -275 -23
rect -255 -45 -251 -43
rect -170 -45 -162 -42
rect -167 -50 -163 -45
rect -79 -48 -71 -45
rect -229 -53 -227 -52
rect -278 -56 -227 -53
rect -296 -80 -292 -77
rect -278 -84 -275 -56
rect -234 -71 -228 -67
rect -242 -84 -239 -81
rect -234 -84 -231 -71
rect -216 -71 -210 -67
rect -76 -53 -72 -48
rect -242 -87 -231 -84
rect -278 -160 -275 -89
rect -234 -96 -231 -87
rect -213 -84 -210 -71
rect -159 -73 -155 -70
rect -204 -77 -166 -73
rect -159 -77 -149 -73
rect -204 -84 -201 -77
rect -159 -82 -155 -77
rect -213 -87 -201 -84
rect -234 -100 -228 -96
rect -213 -96 -210 -87
rect -216 -100 -210 -96
rect -234 -110 -227 -106
rect -258 -132 -250 -129
rect -255 -137 -251 -132
rect -278 -164 -254 -160
rect -247 -161 -243 -157
rect -234 -139 -230 -110
rect -204 -119 -201 -87
rect -152 -87 -149 -77
rect -143 -78 -137 -74
rect -143 -87 -140 -78
rect -125 -78 -119 -74
rect -68 -76 -64 -73
rect -152 -90 -140 -87
rect -197 -99 -191 -95
rect -197 -119 -194 -99
rect -179 -99 -173 -95
rect -204 -122 -194 -119
rect -197 -124 -194 -122
rect -197 -128 -191 -124
rect -176 -122 -173 -99
rect -167 -98 -163 -92
rect -167 -101 -155 -98
rect -159 -107 -155 -101
rect -167 -122 -163 -117
rect -152 -121 -149 -90
rect -143 -103 -140 -90
rect -122 -94 -119 -78
rect -113 -80 -75 -76
rect -68 -80 -58 -76
rect -113 -94 -110 -80
rect -68 -85 -64 -80
rect -143 -107 -137 -103
rect -122 -98 -110 -94
rect -122 -103 -119 -98
rect -125 -107 -119 -103
rect -153 -122 -149 -121
rect -176 -124 -163 -122
rect -179 -126 -163 -124
rect -156 -126 -149 -122
rect -143 -122 -136 -118
rect -113 -122 -110 -98
rect -61 -86 -58 -80
rect -47 -86 -43 25
rect -61 -89 -43 -86
rect -32 -22 -29 25
rect -23 -14 -20 34
rect 103 4 106 50
rect 123 45 128 47
rect 111 34 115 37
rect 45 0 47 4
rect 103 2 113 4
rect 105 0 113 2
rect 110 -3 113 0
rect -13 -10 -7 -7
rect 30 -8 36 -6
rect -13 -13 -11 -10
rect 0 -16 4 -9
rect -18 -19 4 -16
rect 8 -22 12 -9
rect 47 -12 53 -9
rect -32 -25 12 -22
rect -76 -101 -72 -95
rect -76 -104 -64 -101
rect -106 -120 -100 -116
rect -106 -122 -103 -120
rect -179 -128 -173 -126
rect -167 -129 -163 -126
rect -234 -143 -190 -139
rect -234 -161 -230 -143
rect -159 -154 -155 -149
rect -160 -157 -152 -154
rect -143 -155 -139 -122
rect -113 -125 -103 -122
rect -106 -145 -103 -125
rect -68 -110 -64 -104
rect -88 -120 -82 -116
rect -85 -125 -82 -120
rect -76 -125 -72 -120
rect -61 -124 -58 -89
rect -62 -125 -58 -124
rect -85 -129 -72 -125
rect -65 -129 -58 -125
rect -106 -149 -100 -145
rect -85 -145 -82 -129
rect -88 -149 -82 -145
rect -76 -132 -72 -129
rect -32 -144 -29 -25
rect 67 -29 76 -27
rect 131 -29 138 -25
rect -23 -114 -20 -36
rect 45 -69 47 -65
rect 45 -77 48 -75
rect 165 -76 168 6
rect 171 -9 174 50
rect 234 7 236 11
rect 287 6 289 7
rect 225 1 227 5
rect 178 -2 183 0
rect 235 -2 241 -1
rect 189 -9 193 -2
rect 171 -13 193 -9
rect 179 -14 182 -13
rect 197 -73 201 -2
rect 234 -5 241 -2
rect 256 -22 265 -20
rect 214 -66 217 -62
rect 236 -64 240 -62
rect 311 -64 314 77
rect 376 44 379 55
rect 484 52 492 55
rect 487 47 491 52
rect 575 49 583 52
rect 425 44 427 45
rect 376 41 427 44
rect 355 18 362 20
rect 326 17 362 18
rect 326 15 358 17
rect 326 10 329 15
rect 323 7 329 10
rect 376 13 379 41
rect 420 26 426 30
rect 412 13 415 16
rect 420 13 423 26
rect 438 26 444 30
rect 578 44 582 49
rect 412 10 423 13
rect 236 -67 314 -64
rect 376 -63 379 8
rect 420 1 423 10
rect 441 13 444 26
rect 495 24 499 27
rect 450 20 488 24
rect 495 20 505 24
rect 450 13 453 20
rect 495 15 499 20
rect 441 10 453 13
rect 420 -3 426 1
rect 441 1 444 10
rect 438 -3 444 1
rect 420 -13 427 -9
rect 396 -35 404 -32
rect 399 -40 403 -35
rect 376 -67 400 -63
rect 407 -64 411 -60
rect 420 -42 424 -13
rect 450 -22 453 10
rect 502 10 505 20
rect 511 19 517 23
rect 511 10 514 19
rect 529 19 535 23
rect 586 21 590 24
rect 502 7 514 10
rect 457 -2 463 2
rect 457 -22 460 -2
rect 475 -2 481 2
rect 450 -25 460 -22
rect 457 -27 460 -25
rect 457 -31 463 -27
rect 478 -25 481 -2
rect 487 -1 491 5
rect 487 -4 499 -1
rect 495 -10 499 -4
rect 487 -25 491 -20
rect 502 -24 505 7
rect 511 -6 514 7
rect 532 3 535 19
rect 541 17 579 21
rect 586 17 596 21
rect 541 3 544 17
rect 586 12 590 17
rect 511 -10 517 -6
rect 532 -1 544 3
rect 532 -6 535 -1
rect 529 -10 535 -6
rect 501 -25 505 -24
rect 478 -27 491 -25
rect 475 -29 491 -27
rect 498 -29 505 -25
rect 511 -25 518 -21
rect 541 -25 544 -1
rect 593 11 596 17
rect 593 8 607 11
rect 578 -4 582 2
rect 578 -7 590 -4
rect 548 -23 554 -19
rect 548 -25 551 -23
rect 475 -31 481 -29
rect 487 -32 491 -29
rect 420 -46 464 -42
rect 420 -64 424 -46
rect 495 -57 499 -52
rect 494 -60 502 -57
rect 511 -58 515 -25
rect 541 -28 551 -25
rect 548 -48 551 -28
rect 586 -13 590 -7
rect 566 -23 572 -19
rect 569 -28 572 -23
rect 578 -28 582 -23
rect 593 -27 596 8
rect 592 -28 596 -27
rect 569 -32 582 -28
rect 589 -32 596 -28
rect 548 -52 554 -48
rect 569 -48 572 -32
rect 566 -52 572 -48
rect 578 -35 582 -32
rect 511 -62 555 -58
rect 586 -60 590 -55
rect 511 -64 516 -62
rect 585 -63 593 -60
rect 407 -65 412 -64
rect 420 -65 516 -64
rect 236 -73 240 -67
rect 197 -76 240 -73
rect 78 -80 94 -76
rect 111 -80 168 -76
rect 78 -108 81 -80
rect 89 -87 91 -83
rect 76 -112 81 -108
rect -23 -117 24 -114
rect 51 -142 57 -139
rect 29 -144 35 -142
rect -32 -147 35 -144
rect -143 -159 -99 -155
rect -68 -157 -64 -152
rect -143 -161 -138 -159
rect -69 -160 -61 -157
rect -247 -162 -242 -161
rect -234 -162 -138 -161
rect -278 -187 -275 -164
rect -247 -165 -138 -162
rect 78 -162 81 -112
rect 131 -116 281 -113
rect 105 -142 108 -139
rect -247 -169 -243 -165
rect 78 -166 202 -162
rect -255 -184 -251 -179
rect -279 -194 -275 -187
rect 171 -188 232 -184
rect -171 -191 -163 -188
rect -279 -199 -276 -194
rect -168 -196 -164 -191
rect -80 -194 -72 -191
rect -230 -199 -228 -198
rect -279 -202 -228 -199
rect -297 -225 -293 -222
rect -279 -230 -276 -202
rect -235 -217 -229 -213
rect -243 -230 -240 -226
rect -235 -230 -232 -217
rect -217 -217 -211 -213
rect -77 -199 -73 -194
rect 14 -195 75 -191
rect 171 -193 175 -188
rect -243 -233 -232 -230
rect -279 -306 -276 -235
rect -235 -242 -232 -233
rect -214 -230 -211 -217
rect -160 -219 -156 -216
rect -205 -223 -167 -219
rect -160 -223 -150 -219
rect -205 -230 -202 -223
rect -160 -228 -156 -223
rect -214 -233 -202 -230
rect -235 -246 -229 -242
rect -214 -242 -211 -233
rect -217 -246 -211 -242
rect -235 -256 -228 -252
rect -259 -278 -251 -275
rect -256 -283 -252 -278
rect -279 -310 -255 -306
rect -248 -307 -244 -303
rect -235 -285 -231 -256
rect -205 -265 -202 -233
rect -153 -233 -150 -223
rect -144 -224 -138 -220
rect -144 -233 -141 -224
rect 14 -200 18 -195
rect -12 -204 18 -200
rect -8 -208 -4 -204
rect 14 -208 18 -204
rect -126 -224 -120 -220
rect -69 -222 -65 -219
rect -53 -215 -21 -212
rect -153 -236 -141 -233
rect -198 -245 -192 -241
rect -198 -265 -195 -245
rect -180 -245 -174 -241
rect -205 -268 -195 -265
rect -198 -270 -195 -268
rect -198 -274 -192 -270
rect -177 -268 -174 -245
rect -168 -244 -164 -238
rect -168 -247 -156 -244
rect -160 -253 -156 -247
rect -168 -268 -164 -263
rect -153 -267 -150 -236
rect -144 -249 -141 -236
rect -123 -240 -120 -224
rect -114 -226 -76 -222
rect -69 -226 -59 -222
rect -114 -240 -111 -226
rect -69 -231 -65 -226
rect -144 -253 -138 -249
rect -123 -244 -111 -240
rect -123 -249 -120 -244
rect -126 -253 -120 -249
rect -154 -268 -150 -267
rect -177 -270 -164 -268
rect -180 -272 -164 -270
rect -157 -272 -150 -268
rect -144 -268 -137 -264
rect -114 -268 -111 -244
rect -62 -232 -59 -226
rect -53 -232 -50 -215
rect -62 -235 -50 -232
rect -44 -224 -30 -221
rect -77 -247 -73 -241
rect -77 -250 -65 -247
rect -107 -266 -101 -262
rect -107 -268 -104 -266
rect -180 -274 -174 -272
rect -168 -275 -164 -272
rect -235 -289 -191 -285
rect -235 -307 -231 -289
rect -160 -300 -156 -295
rect -161 -303 -153 -300
rect -144 -301 -140 -268
rect -114 -271 -104 -268
rect -107 -291 -104 -271
rect -69 -256 -65 -250
rect -89 -266 -83 -262
rect -86 -271 -83 -266
rect -77 -271 -73 -266
rect -62 -270 -59 -235
rect -44 -259 -41 -224
rect -63 -271 -59 -270
rect -86 -275 -73 -271
rect -66 -275 -59 -271
rect -48 -262 -41 -259
rect -107 -295 -101 -291
rect -86 -291 -83 -275
rect -89 -295 -83 -291
rect -77 -278 -73 -275
rect -144 -305 -100 -301
rect -69 -303 -65 -298
rect -144 -307 -139 -305
rect -70 -306 -62 -303
rect -248 -308 -243 -307
rect -235 -308 -139 -307
rect -279 -340 -276 -310
rect -248 -311 -139 -308
rect -248 -315 -244 -311
rect -256 -330 -252 -325
rect -171 -332 -163 -329
rect -168 -337 -164 -332
rect -80 -335 -72 -332
rect -230 -340 -228 -339
rect -279 -343 -228 -340
rect -297 -367 -293 -364
rect -279 -371 -276 -343
rect -235 -358 -229 -354
rect -243 -371 -240 -368
rect -235 -371 -232 -358
rect -217 -358 -211 -354
rect -77 -340 -73 -335
rect -243 -374 -232 -371
rect -279 -447 -276 -376
rect -235 -383 -232 -374
rect -214 -371 -211 -358
rect -160 -360 -156 -357
rect -205 -364 -167 -360
rect -160 -364 -150 -360
rect -205 -371 -202 -364
rect -160 -369 -156 -364
rect -214 -374 -202 -371
rect -235 -387 -229 -383
rect -214 -383 -211 -374
rect -217 -387 -211 -383
rect -235 -397 -228 -393
rect -259 -419 -251 -416
rect -256 -424 -252 -419
rect -279 -451 -255 -447
rect -248 -448 -244 -444
rect -235 -426 -231 -397
rect -205 -406 -202 -374
rect -153 -374 -150 -364
rect -144 -365 -138 -361
rect -144 -374 -141 -365
rect -126 -365 -120 -361
rect -69 -363 -65 -360
rect -153 -377 -141 -374
rect -198 -386 -192 -382
rect -198 -406 -195 -386
rect -180 -386 -174 -382
rect -205 -409 -195 -406
rect -198 -411 -195 -409
rect -198 -415 -192 -411
rect -177 -409 -174 -386
rect -168 -385 -164 -379
rect -168 -388 -156 -385
rect -160 -394 -156 -388
rect -168 -409 -164 -404
rect -153 -408 -150 -377
rect -144 -390 -141 -377
rect -123 -381 -120 -365
rect -114 -367 -76 -363
rect -69 -367 -59 -363
rect -114 -381 -111 -367
rect -69 -372 -65 -367
rect -144 -394 -138 -390
rect -123 -385 -111 -381
rect -123 -390 -120 -385
rect -126 -394 -120 -390
rect -154 -409 -150 -408
rect -177 -411 -164 -409
rect -180 -413 -164 -411
rect -157 -413 -150 -409
rect -144 -409 -137 -405
rect -114 -409 -111 -385
rect -62 -373 -59 -367
rect -48 -373 -44 -262
rect -62 -376 -44 -373
rect -33 -271 -30 -224
rect -24 -263 -21 -215
rect 31 -199 35 -195
rect 53 -199 57 -195
rect 71 -214 75 -195
rect 149 -197 175 -193
rect 149 -201 153 -197
rect 171 -201 175 -197
rect 71 -218 97 -214
rect 42 -222 46 -219
rect 71 -222 75 -218
rect 93 -222 97 -218
rect 188 -192 192 -188
rect 210 -192 214 -188
rect 228 -207 232 -188
rect 228 -211 254 -207
rect 199 -215 203 -212
rect 228 -215 232 -211
rect 250 -215 254 -211
rect 199 -219 221 -215
rect 42 -226 64 -222
rect 3 -231 7 -228
rect 22 -230 32 -226
rect 22 -231 26 -230
rect 3 -235 26 -231
rect 53 -234 57 -226
rect 14 -243 18 -235
rect -8 -258 -4 -253
rect -12 -262 -4 -258
rect -1 -265 3 -258
rect -19 -268 3 -265
rect 7 -271 11 -258
rect -33 -274 11 -271
rect -77 -388 -73 -382
rect -77 -391 -65 -388
rect -107 -407 -101 -403
rect -107 -409 -104 -407
rect -180 -415 -174 -413
rect -168 -416 -164 -413
rect -235 -430 -191 -426
rect -235 -448 -231 -430
rect -160 -441 -156 -436
rect -161 -444 -153 -441
rect -144 -442 -140 -409
rect -114 -412 -104 -409
rect -107 -432 -104 -412
rect -69 -397 -65 -391
rect -89 -407 -83 -403
rect -86 -412 -83 -407
rect -77 -412 -73 -407
rect -62 -411 -59 -376
rect -33 -393 -30 -274
rect -24 -363 -21 -285
rect 22 -293 26 -235
rect 31 -249 35 -244
rect 44 -249 46 -245
rect 60 -247 64 -226
rect 160 -224 164 -221
rect 179 -223 189 -219
rect 179 -224 183 -223
rect 160 -228 183 -224
rect 210 -227 214 -219
rect 171 -236 175 -228
rect 82 -245 86 -242
rect 29 -255 35 -249
rect 60 -251 72 -247
rect 82 -249 141 -245
rect 81 -256 86 -252
rect 42 -260 46 -257
rect 31 -264 57 -260
rect 31 -268 35 -264
rect 53 -268 57 -264
rect 71 -272 75 -267
rect 66 -276 75 -272
rect 42 -291 46 -288
rect 81 -291 85 -256
rect 93 -257 97 -249
rect 22 -297 32 -293
rect 42 -295 85 -291
rect 53 -303 57 -295
rect 31 -318 35 -313
rect 44 -318 46 -314
rect 26 -322 35 -318
rect 24 -329 60 -326
rect 24 -330 50 -329
rect 24 -334 28 -330
rect 46 -334 50 -330
rect 56 -334 60 -329
rect 35 -357 39 -354
rect 68 -357 72 -354
rect 35 -361 59 -357
rect 68 -361 96 -357
rect 23 -363 25 -362
rect -24 -366 25 -363
rect 46 -369 50 -361
rect 68 -369 72 -361
rect 24 -384 28 -379
rect 22 -385 28 -384
rect 56 -385 60 -379
rect 22 -388 60 -385
rect 28 -393 34 -391
rect -33 -396 34 -393
rect -63 -412 -59 -411
rect -86 -416 -73 -412
rect -66 -416 -59 -412
rect -107 -436 -101 -432
rect -86 -432 -83 -416
rect -89 -436 -83 -432
rect -77 -419 -73 -416
rect 92 -430 96 -361
rect 131 -386 134 -249
rect 138 -258 141 -249
rect 149 -251 153 -246
rect 145 -255 153 -251
rect 156 -258 160 -251
rect 138 -262 160 -258
rect 164 -322 167 -251
rect 179 -286 183 -228
rect 188 -242 192 -237
rect 201 -242 203 -238
rect 217 -240 221 -219
rect 239 -238 243 -235
rect 186 -248 192 -242
rect 217 -244 229 -240
rect 239 -242 256 -238
rect 250 -243 256 -242
rect 238 -249 243 -245
rect 199 -253 203 -250
rect 188 -257 214 -253
rect 188 -261 192 -257
rect 210 -261 214 -257
rect 228 -265 232 -260
rect 223 -269 232 -265
rect 199 -284 203 -281
rect 238 -284 242 -249
rect 250 -250 254 -243
rect 179 -290 189 -286
rect 199 -288 242 -284
rect 210 -296 214 -288
rect 188 -311 192 -306
rect 183 -315 192 -311
rect 203 -313 207 -311
rect 278 -313 281 -116
rect 303 -165 372 -162
rect 203 -316 281 -313
rect 203 -322 206 -316
rect 164 -325 206 -322
rect 369 -338 372 -165
rect 149 -341 372 -338
rect 376 -216 379 -67
rect 407 -68 516 -65
rect 407 -72 411 -68
rect 399 -87 403 -82
rect 484 -208 492 -205
rect 487 -213 491 -208
rect 575 -211 583 -208
rect 425 -216 427 -215
rect 376 -219 427 -216
rect 376 -247 379 -219
rect 420 -234 426 -230
rect 412 -247 415 -244
rect 420 -247 423 -234
rect 438 -234 444 -230
rect 578 -216 582 -211
rect 412 -250 423 -247
rect 376 -323 379 -252
rect 420 -259 423 -250
rect 441 -247 444 -234
rect 495 -236 499 -233
rect 450 -240 488 -236
rect 495 -240 505 -236
rect 450 -247 453 -240
rect 495 -245 499 -240
rect 441 -250 453 -247
rect 420 -263 426 -259
rect 441 -259 444 -250
rect 438 -263 444 -259
rect 420 -273 427 -269
rect 396 -295 404 -292
rect 399 -300 403 -295
rect 376 -327 400 -323
rect 407 -324 411 -320
rect 420 -302 424 -273
rect 450 -282 453 -250
rect 502 -250 505 -240
rect 511 -241 517 -237
rect 511 -250 514 -241
rect 529 -241 535 -237
rect 586 -239 590 -236
rect 502 -253 514 -250
rect 457 -262 463 -258
rect 457 -282 460 -262
rect 475 -262 481 -258
rect 450 -285 460 -282
rect 457 -287 460 -285
rect 457 -291 463 -287
rect 478 -285 481 -262
rect 487 -261 491 -255
rect 487 -264 499 -261
rect 495 -270 499 -264
rect 487 -285 491 -280
rect 502 -284 505 -253
rect 511 -266 514 -253
rect 532 -257 535 -241
rect 541 -243 579 -239
rect 586 -243 596 -239
rect 541 -257 544 -243
rect 586 -248 590 -243
rect 511 -270 517 -266
rect 532 -261 544 -257
rect 532 -266 535 -261
rect 529 -270 535 -266
rect 501 -285 505 -284
rect 478 -287 491 -285
rect 475 -289 491 -287
rect 498 -289 505 -285
rect 511 -285 518 -281
rect 541 -285 544 -261
rect 593 -249 596 -243
rect 593 -252 607 -249
rect 578 -264 582 -258
rect 578 -267 590 -264
rect 548 -283 554 -279
rect 548 -285 551 -283
rect 475 -291 481 -289
rect 487 -292 491 -289
rect 420 -306 464 -302
rect 420 -324 424 -306
rect 495 -317 499 -312
rect 494 -320 502 -317
rect 511 -318 515 -285
rect 541 -288 551 -285
rect 548 -308 551 -288
rect 586 -273 590 -267
rect 566 -283 572 -279
rect 569 -288 572 -283
rect 578 -288 582 -283
rect 593 -287 596 -252
rect 592 -288 596 -287
rect 569 -292 582 -288
rect 589 -292 596 -288
rect 548 -312 554 -308
rect 569 -308 572 -292
rect 566 -312 572 -308
rect 578 -295 582 -292
rect 511 -322 555 -318
rect 586 -320 590 -315
rect 511 -324 516 -322
rect 585 -323 593 -320
rect 407 -325 412 -324
rect 420 -325 516 -324
rect 149 -342 154 -341
rect 140 -353 176 -350
rect 140 -354 166 -353
rect 140 -358 144 -354
rect 162 -358 166 -354
rect 172 -358 176 -353
rect 191 -353 215 -349
rect 232 -353 269 -349
rect 151 -381 155 -378
rect 184 -381 188 -378
rect 191 -380 194 -353
rect 210 -359 243 -356
rect 210 -360 217 -359
rect 213 -363 217 -360
rect 239 -363 243 -359
rect 151 -385 175 -381
rect 184 -385 191 -381
rect 131 -390 141 -386
rect 154 -392 155 -388
rect 162 -393 166 -385
rect 184 -393 188 -385
rect 230 -386 234 -383
rect 247 -386 251 -383
rect 222 -390 240 -386
rect 247 -389 255 -386
rect 222 -395 226 -390
rect 247 -395 251 -389
rect 140 -409 144 -403
rect 172 -409 176 -403
rect 140 -412 176 -409
rect 213 -409 217 -405
rect 231 -409 235 -405
rect 239 -409 243 -405
rect 213 -412 243 -409
rect 157 -416 164 -412
rect 226 -415 229 -412
rect 266 -430 269 -353
rect 92 -433 362 -430
rect -144 -446 -100 -442
rect -69 -444 -65 -439
rect -144 -448 -139 -446
rect -70 -447 -62 -444
rect -248 -449 -243 -448
rect -235 -449 -139 -448
rect -279 -471 -276 -451
rect -248 -452 -139 -449
rect -248 -456 -244 -452
rect 256 -456 259 -443
rect 256 -459 287 -456
rect -256 -471 -252 -466
rect -280 -478 -276 -471
rect -172 -475 -164 -472
rect 177 -473 238 -469
rect -280 -483 -277 -478
rect -169 -480 -165 -475
rect -81 -478 -73 -475
rect -231 -483 -229 -482
rect -280 -486 -229 -483
rect -298 -509 -294 -506
rect -280 -514 -277 -486
rect -236 -501 -230 -497
rect -244 -514 -241 -510
rect -236 -514 -233 -501
rect -218 -501 -212 -497
rect -78 -483 -74 -478
rect 20 -480 81 -476
rect 177 -478 181 -473
rect -244 -517 -233 -514
rect -280 -582 -277 -519
rect -236 -526 -233 -517
rect -215 -514 -212 -501
rect -161 -503 -157 -500
rect -206 -507 -168 -503
rect -161 -507 -151 -503
rect -206 -514 -203 -507
rect -161 -512 -157 -507
rect -215 -517 -203 -514
rect -236 -530 -230 -526
rect -215 -526 -212 -517
rect -218 -530 -212 -526
rect -236 -540 -229 -536
rect -260 -562 -252 -559
rect -282 -590 -277 -582
rect -257 -567 -253 -562
rect -282 -594 -256 -590
rect -249 -591 -245 -587
rect -236 -569 -232 -540
rect -206 -549 -203 -517
rect -154 -517 -151 -507
rect -145 -508 -139 -504
rect -145 -517 -142 -508
rect 20 -485 24 -480
rect -6 -489 24 -485
rect -2 -493 2 -489
rect 20 -493 24 -489
rect -127 -508 -121 -504
rect -70 -506 -66 -503
rect -54 -500 -15 -497
rect -154 -520 -142 -517
rect -199 -529 -193 -525
rect -199 -549 -196 -529
rect -181 -529 -175 -525
rect -206 -552 -196 -549
rect -199 -554 -196 -552
rect -199 -558 -193 -554
rect -178 -552 -175 -529
rect -169 -528 -165 -522
rect -169 -531 -157 -528
rect -161 -537 -157 -531
rect -169 -552 -165 -547
rect -154 -551 -151 -520
rect -145 -533 -142 -520
rect -124 -524 -121 -508
rect -115 -510 -77 -506
rect -70 -510 -60 -506
rect -115 -524 -112 -510
rect -70 -515 -66 -510
rect -145 -537 -139 -533
rect -124 -528 -112 -524
rect -124 -533 -121 -528
rect -127 -537 -121 -533
rect -155 -552 -151 -551
rect -178 -554 -165 -552
rect -181 -556 -165 -554
rect -158 -556 -151 -552
rect -145 -552 -138 -548
rect -115 -552 -112 -528
rect -63 -516 -60 -510
rect -54 -516 -51 -500
rect -63 -519 -51 -516
rect -45 -509 -24 -506
rect -78 -531 -74 -525
rect -78 -534 -66 -531
rect -108 -550 -102 -546
rect -108 -552 -105 -550
rect -181 -558 -175 -556
rect -169 -559 -165 -556
rect -236 -573 -192 -569
rect -236 -591 -232 -573
rect -161 -584 -157 -579
rect -162 -587 -154 -584
rect -145 -585 -141 -552
rect -115 -555 -105 -552
rect -108 -575 -105 -555
rect -70 -540 -66 -534
rect -90 -550 -84 -546
rect -87 -555 -84 -550
rect -78 -555 -74 -550
rect -63 -554 -60 -519
rect -45 -543 -42 -509
rect -64 -555 -60 -554
rect -87 -559 -74 -555
rect -67 -559 -60 -555
rect -49 -546 -42 -543
rect -108 -579 -102 -575
rect -87 -575 -84 -559
rect -90 -579 -84 -575
rect -78 -562 -74 -559
rect -145 -589 -101 -585
rect -70 -587 -66 -582
rect -145 -591 -140 -589
rect -71 -590 -63 -587
rect -249 -592 -244 -591
rect -236 -592 -140 -591
rect -282 -624 -277 -594
rect -249 -595 -140 -592
rect -249 -599 -245 -595
rect -257 -614 -253 -609
rect -172 -616 -164 -613
rect -169 -621 -165 -616
rect -81 -619 -73 -616
rect -231 -624 -229 -623
rect -282 -627 -229 -624
rect -298 -651 -294 -648
rect -282 -655 -277 -627
rect -236 -642 -230 -638
rect -244 -655 -241 -652
rect -236 -655 -233 -642
rect -218 -642 -212 -638
rect -78 -624 -74 -619
rect -282 -660 -280 -655
rect -244 -658 -233 -655
rect -282 -731 -277 -660
rect -236 -667 -233 -658
rect -215 -655 -212 -642
rect -161 -644 -157 -641
rect -206 -648 -168 -644
rect -161 -648 -151 -644
rect -206 -655 -203 -648
rect -161 -653 -157 -648
rect -215 -658 -203 -655
rect -236 -671 -230 -667
rect -215 -667 -212 -658
rect -218 -671 -212 -667
rect -236 -681 -229 -677
rect -260 -703 -252 -700
rect -257 -708 -253 -703
rect -282 -735 -256 -731
rect -249 -732 -245 -728
rect -236 -710 -232 -681
rect -206 -690 -203 -658
rect -154 -658 -151 -648
rect -145 -649 -139 -645
rect -145 -658 -142 -649
rect -127 -649 -121 -645
rect -70 -647 -66 -644
rect -154 -661 -142 -658
rect -199 -670 -193 -666
rect -199 -690 -196 -670
rect -181 -670 -175 -666
rect -206 -693 -196 -690
rect -199 -695 -196 -693
rect -199 -699 -193 -695
rect -178 -693 -175 -670
rect -169 -669 -165 -663
rect -169 -672 -157 -669
rect -161 -678 -157 -672
rect -169 -693 -165 -688
rect -154 -692 -151 -661
rect -145 -674 -142 -661
rect -124 -665 -121 -649
rect -115 -651 -77 -647
rect -70 -651 -60 -647
rect -115 -665 -112 -651
rect -70 -656 -66 -651
rect -145 -678 -139 -674
rect -124 -669 -112 -665
rect -124 -674 -121 -669
rect -127 -678 -121 -674
rect -155 -693 -151 -692
rect -178 -695 -165 -693
rect -181 -697 -165 -695
rect -158 -697 -151 -693
rect -145 -693 -138 -689
rect -115 -693 -112 -669
rect -63 -657 -60 -651
rect -49 -657 -45 -546
rect -63 -660 -45 -657
rect -27 -556 -24 -509
rect -18 -548 -15 -500
rect 37 -484 41 -480
rect 59 -484 63 -480
rect 77 -499 81 -480
rect 155 -482 181 -478
rect 155 -486 159 -482
rect 177 -486 181 -482
rect 77 -503 103 -499
rect 48 -507 52 -504
rect 77 -507 81 -503
rect 99 -507 103 -503
rect 194 -477 198 -473
rect 216 -477 220 -473
rect 234 -492 238 -473
rect 234 -496 260 -492
rect 205 -500 209 -497
rect 234 -500 238 -496
rect 256 -500 260 -496
rect 205 -504 227 -500
rect 48 -511 70 -507
rect 9 -516 13 -513
rect 28 -515 38 -511
rect 28 -516 32 -515
rect 9 -520 32 -516
rect 59 -519 63 -511
rect 20 -528 24 -520
rect -2 -543 2 -538
rect -6 -547 2 -543
rect 5 -550 9 -543
rect -13 -553 9 -550
rect 13 -556 17 -543
rect -27 -559 17 -556
rect -78 -672 -74 -666
rect -78 -675 -66 -672
rect -108 -691 -102 -687
rect -108 -693 -105 -691
rect -181 -699 -175 -697
rect -169 -700 -165 -697
rect -236 -714 -192 -710
rect -236 -732 -232 -714
rect -161 -725 -157 -720
rect -162 -728 -154 -725
rect -145 -726 -141 -693
rect -115 -696 -105 -693
rect -108 -716 -105 -696
rect -70 -681 -66 -675
rect -90 -691 -84 -687
rect -87 -696 -84 -691
rect -78 -696 -74 -691
rect -63 -695 -60 -660
rect -27 -678 -24 -559
rect -18 -648 -15 -570
rect 28 -578 32 -520
rect 37 -534 41 -529
rect 50 -534 52 -530
rect 66 -532 70 -511
rect 166 -509 170 -506
rect 185 -508 195 -504
rect 185 -509 189 -508
rect 166 -513 189 -509
rect 216 -512 220 -504
rect 177 -521 181 -513
rect 88 -530 92 -527
rect 35 -540 41 -534
rect 66 -536 78 -532
rect 88 -534 147 -530
rect 87 -541 92 -537
rect 48 -545 52 -542
rect 37 -549 63 -545
rect 37 -553 41 -549
rect 59 -553 63 -549
rect 77 -557 81 -552
rect 72 -561 81 -557
rect 48 -576 52 -573
rect 87 -576 91 -541
rect 99 -542 103 -534
rect 28 -582 38 -578
rect 48 -580 91 -576
rect 59 -588 63 -580
rect 37 -603 41 -598
rect 50 -603 52 -599
rect 32 -607 41 -603
rect 30 -614 66 -611
rect 30 -615 56 -614
rect 30 -619 34 -615
rect 52 -619 56 -615
rect 62 -619 66 -614
rect 41 -642 45 -639
rect 74 -642 78 -639
rect 41 -646 65 -642
rect 74 -646 89 -642
rect 29 -648 31 -647
rect -18 -651 31 -648
rect 52 -654 56 -646
rect 74 -654 78 -646
rect 30 -669 34 -664
rect 28 -670 34 -669
rect 62 -670 66 -664
rect 28 -673 66 -670
rect 34 -678 40 -676
rect -27 -681 40 -678
rect -64 -696 -60 -695
rect -87 -700 -74 -696
rect -67 -700 -60 -696
rect -108 -720 -102 -716
rect -87 -716 -84 -700
rect -90 -720 -84 -716
rect -78 -703 -74 -700
rect -145 -730 -101 -726
rect -70 -728 -66 -723
rect -145 -732 -140 -730
rect -71 -731 -63 -728
rect -249 -733 -244 -732
rect -236 -733 -140 -732
rect -282 -772 -277 -735
rect -249 -736 -140 -733
rect -249 -740 -245 -736
rect -257 -755 -253 -750
rect -172 -764 -164 -762
rect -169 -769 -165 -764
rect -81 -767 -73 -764
rect -231 -772 -229 -771
rect -282 -775 -229 -772
rect -298 -798 -294 -795
rect -282 -803 -277 -775
rect -236 -790 -230 -786
rect -244 -803 -241 -799
rect -236 -803 -233 -790
rect -218 -790 -212 -786
rect -78 -772 -74 -767
rect -282 -808 -280 -803
rect -244 -806 -233 -803
rect -282 -879 -277 -808
rect -236 -815 -233 -806
rect -215 -803 -212 -790
rect -161 -792 -157 -789
rect -206 -796 -168 -792
rect -161 -796 -151 -792
rect -206 -803 -203 -796
rect -161 -801 -157 -796
rect -215 -806 -203 -803
rect -236 -819 -230 -815
rect -215 -815 -212 -806
rect -218 -819 -212 -815
rect -236 -829 -229 -825
rect -260 -851 -252 -848
rect -257 -856 -253 -851
rect -282 -883 -256 -879
rect -249 -880 -245 -876
rect -236 -858 -232 -829
rect -206 -838 -203 -806
rect -154 -806 -151 -796
rect -145 -797 -139 -793
rect -145 -806 -142 -797
rect -127 -797 -121 -793
rect -70 -795 -66 -792
rect -154 -809 -142 -806
rect -199 -818 -193 -814
rect -199 -838 -196 -818
rect -181 -818 -175 -814
rect -206 -841 -196 -838
rect -199 -843 -196 -841
rect -199 -847 -193 -843
rect -178 -841 -175 -818
rect -169 -817 -165 -811
rect -169 -820 -157 -817
rect -161 -826 -157 -820
rect -169 -841 -165 -836
rect -154 -840 -151 -809
rect -145 -822 -142 -809
rect -124 -813 -121 -797
rect -115 -799 -77 -795
rect -70 -799 -60 -795
rect 85 -796 89 -646
rect 137 -671 140 -534
rect 144 -543 147 -534
rect 155 -536 159 -531
rect 151 -540 159 -536
rect 162 -543 166 -536
rect 144 -547 166 -543
rect 170 -607 173 -536
rect 185 -571 189 -513
rect 194 -527 198 -522
rect 207 -527 209 -523
rect 223 -525 227 -504
rect 245 -523 249 -520
rect 192 -533 198 -527
rect 223 -529 235 -525
rect 245 -527 262 -523
rect 256 -528 262 -527
rect 244 -534 249 -530
rect 205 -538 209 -535
rect 194 -542 220 -538
rect 194 -546 198 -542
rect 216 -546 220 -542
rect 234 -550 238 -545
rect 229 -554 238 -550
rect 205 -569 209 -566
rect 244 -569 248 -534
rect 256 -535 260 -528
rect 185 -575 195 -571
rect 205 -573 248 -569
rect 216 -581 220 -573
rect 194 -596 198 -591
rect 189 -600 198 -596
rect 209 -598 213 -596
rect 284 -598 287 -459
rect 209 -601 287 -598
rect 209 -607 212 -601
rect 170 -610 212 -607
rect 359 -621 362 -433
rect 155 -624 362 -621
rect 376 -500 379 -327
rect 407 -328 516 -325
rect 407 -332 411 -328
rect 399 -347 403 -342
rect 484 -492 492 -489
rect 487 -497 491 -492
rect 575 -495 583 -492
rect 425 -500 427 -499
rect 376 -503 427 -500
rect 376 -531 379 -503
rect 420 -518 426 -514
rect 412 -531 415 -528
rect 420 -531 423 -518
rect 438 -518 444 -514
rect 578 -500 582 -495
rect 412 -534 423 -531
rect 376 -607 379 -536
rect 420 -543 423 -534
rect 441 -531 444 -518
rect 495 -520 499 -517
rect 450 -524 488 -520
rect 495 -524 505 -520
rect 450 -531 453 -524
rect 495 -529 499 -524
rect 441 -534 453 -531
rect 420 -547 426 -543
rect 441 -543 444 -534
rect 438 -547 444 -543
rect 420 -557 427 -553
rect 396 -579 404 -576
rect 399 -584 403 -579
rect 376 -611 400 -607
rect 407 -608 411 -604
rect 420 -586 424 -557
rect 450 -566 453 -534
rect 502 -534 505 -524
rect 511 -525 517 -521
rect 511 -534 514 -525
rect 529 -525 535 -521
rect 586 -523 590 -520
rect 502 -537 514 -534
rect 457 -546 463 -542
rect 457 -566 460 -546
rect 475 -546 481 -542
rect 450 -569 460 -566
rect 457 -571 460 -569
rect 457 -575 463 -571
rect 478 -569 481 -546
rect 487 -545 491 -539
rect 487 -548 499 -545
rect 495 -554 499 -548
rect 487 -569 491 -564
rect 502 -568 505 -537
rect 511 -550 514 -537
rect 532 -541 535 -525
rect 541 -527 579 -523
rect 586 -527 596 -523
rect 541 -541 544 -527
rect 586 -532 590 -527
rect 511 -554 517 -550
rect 532 -545 544 -541
rect 532 -550 535 -545
rect 529 -554 535 -550
rect 501 -569 505 -568
rect 478 -571 491 -569
rect 475 -573 491 -571
rect 498 -573 505 -569
rect 511 -569 518 -565
rect 541 -569 544 -545
rect 593 -533 596 -527
rect 593 -536 607 -533
rect 578 -548 582 -542
rect 578 -551 590 -548
rect 548 -567 554 -563
rect 548 -569 551 -567
rect 475 -575 481 -573
rect 487 -576 491 -573
rect 420 -590 464 -586
rect 420 -608 424 -590
rect 495 -601 499 -596
rect 494 -604 502 -601
rect 511 -602 515 -569
rect 541 -572 551 -569
rect 548 -592 551 -572
rect 586 -557 590 -551
rect 566 -567 572 -563
rect 569 -572 572 -567
rect 578 -572 582 -567
rect 593 -571 596 -536
rect 592 -572 596 -571
rect 569 -576 582 -572
rect 589 -576 596 -572
rect 548 -596 554 -592
rect 569 -592 572 -576
rect 566 -596 572 -592
rect 578 -579 582 -576
rect 511 -606 555 -602
rect 586 -604 590 -599
rect 511 -608 516 -606
rect 585 -607 593 -604
rect 407 -609 412 -608
rect 420 -609 516 -608
rect 155 -627 160 -624
rect 207 -631 308 -628
rect 207 -634 211 -631
rect 304 -634 308 -631
rect 146 -638 182 -635
rect 146 -639 172 -638
rect 146 -643 150 -639
rect 168 -643 172 -639
rect 178 -643 182 -638
rect 197 -638 211 -634
rect 219 -638 255 -635
rect 157 -666 161 -663
rect 190 -666 194 -663
rect 197 -664 200 -638
rect 219 -639 245 -638
rect 219 -643 223 -639
rect 241 -643 245 -639
rect 251 -643 255 -638
rect 270 -638 291 -634
rect 157 -670 181 -666
rect 190 -670 197 -666
rect 230 -666 234 -663
rect 263 -666 267 -663
rect 270 -665 273 -638
rect 286 -644 319 -641
rect 286 -645 293 -644
rect 289 -648 293 -645
rect 315 -648 319 -644
rect 230 -670 254 -666
rect 263 -670 270 -666
rect 137 -675 147 -671
rect 137 -704 140 -675
rect 160 -677 161 -673
rect 168 -678 172 -670
rect 190 -678 194 -670
rect 213 -675 220 -671
rect 146 -694 150 -688
rect 178 -694 182 -688
rect 146 -697 182 -694
rect 163 -701 170 -697
rect 213 -704 216 -675
rect 233 -677 234 -673
rect 241 -678 245 -670
rect 263 -678 267 -670
rect 306 -671 310 -668
rect 323 -671 327 -668
rect 298 -675 316 -671
rect 323 -674 334 -671
rect 298 -680 302 -675
rect 323 -680 327 -674
rect 219 -694 223 -688
rect 251 -694 255 -688
rect 219 -697 255 -694
rect 289 -694 293 -690
rect 307 -694 311 -690
rect 315 -694 319 -690
rect 289 -697 319 -694
rect 236 -701 243 -697
rect 302 -700 305 -697
rect 137 -707 216 -704
rect 330 -709 334 -674
rect 244 -712 334 -709
rect 244 -715 248 -712
rect 261 -719 298 -715
rect 239 -725 272 -722
rect 239 -726 246 -725
rect 242 -729 246 -726
rect 268 -729 272 -725
rect 259 -752 263 -749
rect 276 -752 280 -749
rect 251 -756 269 -752
rect 276 -755 284 -752
rect 251 -761 255 -756
rect 276 -761 280 -755
rect 242 -775 246 -771
rect 260 -775 264 -771
rect 268 -775 272 -771
rect 242 -778 272 -775
rect 255 -781 258 -778
rect 295 -796 298 -719
rect 376 -769 379 -611
rect 407 -612 516 -609
rect 407 -616 411 -612
rect 399 -631 403 -626
rect 484 -761 492 -758
rect 487 -766 491 -761
rect 575 -764 583 -761
rect 425 -769 427 -768
rect 376 -772 427 -769
rect 85 -799 352 -796
rect -115 -813 -112 -799
rect -70 -804 -66 -799
rect -145 -826 -139 -822
rect -124 -817 -112 -813
rect -124 -822 -121 -817
rect -127 -826 -121 -822
rect -155 -841 -151 -840
rect -178 -843 -165 -841
rect -181 -845 -165 -843
rect -158 -845 -151 -841
rect -145 -841 -138 -837
rect -115 -841 -112 -817
rect -63 -805 -60 -799
rect -63 -808 -51 -805
rect -78 -820 -74 -814
rect -78 -823 -66 -820
rect -108 -839 -102 -835
rect -108 -841 -105 -839
rect -181 -847 -175 -845
rect -169 -848 -165 -845
rect -236 -862 -192 -858
rect -236 -880 -232 -862
rect -161 -873 -157 -868
rect -162 -876 -154 -873
rect -145 -874 -141 -841
rect -115 -844 -105 -841
rect -108 -864 -105 -844
rect -70 -829 -66 -823
rect -90 -839 -84 -835
rect -87 -844 -84 -839
rect -78 -844 -74 -839
rect -63 -843 -60 -808
rect -64 -844 -60 -843
rect -87 -848 -74 -844
rect -67 -848 -60 -844
rect -108 -868 -102 -864
rect -87 -864 -84 -848
rect -90 -868 -84 -864
rect -78 -851 -74 -848
rect -145 -878 -101 -874
rect -70 -876 -66 -871
rect -145 -880 -140 -878
rect -71 -879 -63 -876
rect -54 -877 -51 -808
rect 285 -837 288 -809
rect 284 -840 288 -837
rect 177 -853 238 -849
rect 20 -860 81 -856
rect 177 -858 181 -853
rect 20 -865 24 -860
rect -6 -869 24 -865
rect -2 -873 2 -869
rect 20 -873 24 -869
rect -54 -880 -15 -877
rect -249 -881 -244 -880
rect -236 -881 -140 -880
rect -282 -913 -277 -883
rect -249 -884 -140 -881
rect -249 -888 -245 -884
rect -49 -889 -24 -886
rect -257 -903 -253 -898
rect -172 -905 -164 -902
rect -169 -910 -165 -905
rect -81 -908 -73 -905
rect -231 -913 -229 -912
rect -282 -916 -229 -913
rect -298 -940 -294 -937
rect -282 -944 -277 -916
rect -236 -931 -230 -927
rect -244 -944 -241 -941
rect -236 -944 -233 -931
rect -218 -931 -212 -927
rect -78 -913 -74 -908
rect -282 -949 -280 -944
rect -244 -947 -233 -944
rect -282 -1020 -277 -949
rect -236 -956 -233 -947
rect -215 -944 -212 -931
rect -161 -933 -157 -930
rect -206 -937 -168 -933
rect -161 -937 -151 -933
rect -206 -944 -203 -937
rect -161 -942 -157 -937
rect -215 -947 -203 -944
rect -236 -960 -230 -956
rect -215 -956 -212 -947
rect -218 -960 -212 -956
rect -236 -970 -229 -966
rect -260 -992 -252 -989
rect -257 -997 -253 -992
rect -282 -1024 -256 -1020
rect -249 -1021 -245 -1017
rect -236 -999 -232 -970
rect -206 -979 -203 -947
rect -154 -947 -151 -937
rect -145 -938 -139 -934
rect -145 -947 -142 -938
rect -127 -938 -121 -934
rect -70 -936 -66 -933
rect -154 -950 -142 -947
rect -199 -959 -193 -955
rect -199 -979 -196 -959
rect -181 -959 -175 -955
rect -206 -982 -196 -979
rect -199 -984 -196 -982
rect -199 -988 -193 -984
rect -178 -982 -175 -959
rect -169 -958 -165 -952
rect -169 -961 -157 -958
rect -161 -967 -157 -961
rect -169 -982 -165 -977
rect -154 -981 -151 -950
rect -145 -963 -142 -950
rect -124 -954 -121 -938
rect -115 -940 -77 -936
rect -70 -940 -60 -936
rect -115 -954 -112 -940
rect -70 -945 -66 -940
rect -145 -967 -139 -963
rect -124 -958 -112 -954
rect -124 -963 -121 -958
rect -127 -967 -121 -963
rect -155 -982 -151 -981
rect -178 -984 -165 -982
rect -181 -986 -165 -984
rect -158 -986 -151 -982
rect -145 -982 -138 -978
rect -115 -982 -112 -958
rect -63 -946 -60 -940
rect -49 -946 -45 -889
rect -63 -949 -45 -946
rect -27 -936 -24 -889
rect -18 -910 -15 -880
rect 37 -864 41 -860
rect 59 -864 63 -860
rect 77 -879 81 -860
rect 155 -862 181 -858
rect 155 -866 159 -862
rect 177 -866 181 -862
rect 77 -883 103 -879
rect 48 -887 52 -884
rect 77 -887 81 -883
rect 99 -887 103 -883
rect 194 -857 198 -853
rect 216 -857 220 -853
rect 234 -872 238 -853
rect 234 -876 260 -872
rect 205 -880 209 -877
rect 234 -880 238 -876
rect 256 -880 260 -876
rect 205 -884 227 -880
rect 48 -891 70 -887
rect 9 -896 13 -893
rect 28 -895 38 -891
rect 28 -896 32 -895
rect 9 -900 32 -896
rect 59 -899 63 -891
rect 20 -908 24 -900
rect -18 -928 -15 -915
rect -2 -923 2 -918
rect -6 -927 2 -923
rect 5 -930 9 -923
rect -13 -933 9 -930
rect 13 -936 17 -923
rect -27 -939 17 -936
rect -78 -961 -74 -955
rect -78 -964 -66 -961
rect -108 -980 -102 -976
rect -108 -982 -105 -980
rect -181 -988 -175 -986
rect -169 -989 -165 -986
rect -236 -1003 -192 -999
rect -236 -1021 -232 -1003
rect -161 -1014 -157 -1009
rect -162 -1017 -154 -1014
rect -145 -1015 -141 -982
rect -115 -985 -105 -982
rect -108 -1005 -105 -985
rect -70 -970 -66 -964
rect -90 -980 -84 -976
rect -87 -985 -84 -980
rect -78 -985 -74 -980
rect -63 -984 -60 -949
rect -27 -979 -24 -939
rect -64 -985 -60 -984
rect -87 -989 -74 -985
rect -67 -989 -60 -985
rect -108 -1009 -102 -1005
rect -87 -1005 -84 -989
rect -90 -1009 -84 -1005
rect -78 -992 -74 -989
rect -145 -1019 -101 -1015
rect -70 -1017 -66 -1012
rect -145 -1021 -140 -1019
rect -71 -1020 -63 -1017
rect -249 -1022 -244 -1021
rect -236 -1022 -140 -1021
rect -282 -1054 -277 -1024
rect -249 -1025 -140 -1022
rect -249 -1029 -245 -1025
rect -257 -1044 -253 -1039
rect -282 -1215 -278 -1054
rect -27 -1058 -24 -984
rect -18 -1028 -15 -950
rect 28 -958 32 -900
rect 37 -914 41 -909
rect 35 -920 41 -914
rect 66 -912 70 -891
rect 166 -889 170 -886
rect 185 -888 195 -884
rect 185 -889 189 -888
rect 166 -893 189 -889
rect 216 -892 220 -884
rect 177 -901 181 -893
rect 88 -910 92 -907
rect 142 -910 147 -908
rect 66 -916 78 -912
rect 88 -914 147 -910
rect 87 -921 92 -917
rect 48 -925 52 -922
rect 37 -929 63 -925
rect 37 -933 41 -929
rect 59 -933 63 -929
rect 77 -937 81 -932
rect 72 -941 81 -937
rect 48 -956 52 -953
rect 87 -956 91 -921
rect 99 -922 103 -914
rect 28 -962 38 -958
rect 48 -960 91 -956
rect 59 -968 63 -960
rect 37 -983 41 -978
rect 32 -987 41 -983
rect 30 -994 66 -991
rect 30 -995 56 -994
rect 30 -999 34 -995
rect 52 -999 56 -995
rect 62 -999 66 -994
rect 41 -1022 45 -1019
rect 74 -1022 78 -1019
rect 41 -1026 65 -1022
rect 74 -1026 89 -1022
rect 29 -1028 31 -1027
rect -18 -1031 31 -1028
rect 52 -1034 56 -1026
rect 74 -1034 78 -1026
rect 30 -1049 34 -1044
rect 28 -1050 34 -1049
rect 62 -1050 66 -1044
rect 28 -1053 66 -1050
rect 34 -1058 40 -1056
rect -27 -1061 40 -1058
rect 85 -1194 89 -1026
rect 137 -1051 140 -914
rect 144 -923 147 -914
rect 155 -916 159 -911
rect 151 -920 159 -916
rect 162 -923 166 -916
rect 144 -927 166 -923
rect 170 -987 173 -916
rect 185 -951 189 -893
rect 194 -907 198 -902
rect 192 -913 198 -907
rect 223 -905 227 -884
rect 245 -903 249 -900
rect 223 -909 235 -905
rect 245 -907 262 -903
rect 256 -908 262 -907
rect 244 -914 249 -910
rect 205 -918 209 -915
rect 194 -922 220 -918
rect 194 -926 198 -922
rect 216 -926 220 -922
rect 234 -930 238 -925
rect 229 -934 238 -930
rect 205 -949 209 -946
rect 244 -949 248 -914
rect 256 -915 260 -908
rect 185 -955 195 -951
rect 205 -953 248 -949
rect 216 -961 220 -953
rect 194 -976 198 -971
rect 189 -980 198 -976
rect 209 -978 213 -976
rect 284 -978 287 -840
rect 296 -907 328 -904
rect 209 -981 287 -978
rect 209 -987 212 -981
rect 170 -990 212 -987
rect 349 -1001 352 -799
rect 155 -1004 352 -1001
rect 376 -800 379 -772
rect 420 -787 426 -783
rect 412 -800 415 -797
rect 420 -800 423 -787
rect 438 -787 444 -783
rect 578 -769 582 -764
rect 412 -803 423 -800
rect 376 -876 379 -805
rect 420 -812 423 -803
rect 441 -800 444 -787
rect 495 -789 499 -786
rect 450 -793 488 -789
rect 495 -793 505 -789
rect 450 -800 453 -793
rect 495 -798 499 -793
rect 441 -803 453 -800
rect 420 -816 426 -812
rect 441 -812 444 -803
rect 438 -816 444 -812
rect 420 -826 427 -822
rect 396 -848 404 -845
rect 399 -853 403 -848
rect 376 -880 400 -876
rect 407 -877 411 -873
rect 420 -855 424 -826
rect 450 -835 453 -803
rect 502 -803 505 -793
rect 511 -794 517 -790
rect 511 -803 514 -794
rect 529 -794 535 -790
rect 586 -792 590 -789
rect 502 -806 514 -803
rect 457 -815 463 -811
rect 457 -835 460 -815
rect 475 -815 481 -811
rect 450 -838 460 -835
rect 457 -840 460 -838
rect 457 -844 463 -840
rect 478 -838 481 -815
rect 487 -814 491 -808
rect 487 -817 499 -814
rect 495 -823 499 -817
rect 487 -838 491 -833
rect 502 -837 505 -806
rect 511 -819 514 -806
rect 532 -810 535 -794
rect 541 -796 579 -792
rect 586 -796 596 -792
rect 541 -810 544 -796
rect 586 -801 590 -796
rect 511 -823 517 -819
rect 532 -814 544 -810
rect 532 -819 535 -814
rect 529 -823 535 -819
rect 501 -838 505 -837
rect 478 -840 491 -838
rect 475 -842 491 -840
rect 498 -842 505 -838
rect 511 -838 518 -834
rect 541 -838 544 -814
rect 593 -802 596 -796
rect 593 -805 607 -802
rect 578 -817 582 -811
rect 578 -820 590 -817
rect 548 -836 554 -832
rect 548 -838 551 -836
rect 475 -844 481 -842
rect 487 -845 491 -842
rect 420 -859 464 -855
rect 420 -877 424 -859
rect 495 -870 499 -865
rect 494 -873 502 -870
rect 511 -871 515 -838
rect 541 -841 551 -838
rect 548 -861 551 -841
rect 586 -826 590 -820
rect 566 -836 572 -832
rect 569 -841 572 -836
rect 578 -841 582 -836
rect 593 -840 596 -805
rect 592 -841 596 -840
rect 569 -845 582 -841
rect 589 -845 596 -841
rect 548 -865 554 -861
rect 569 -861 572 -845
rect 566 -865 572 -861
rect 578 -848 582 -845
rect 511 -875 555 -871
rect 586 -873 590 -868
rect 511 -877 516 -875
rect 585 -876 593 -873
rect 407 -878 412 -877
rect 420 -878 516 -877
rect 376 -988 379 -880
rect 407 -881 516 -878
rect 407 -885 411 -881
rect 399 -900 403 -895
rect 484 -980 492 -977
rect 487 -985 491 -980
rect 575 -983 583 -980
rect 425 -988 427 -987
rect 376 -991 427 -988
rect 155 -1007 160 -1004
rect 207 -1011 309 -1008
rect 207 -1014 211 -1011
rect 305 -1014 309 -1011
rect 146 -1018 182 -1015
rect 146 -1019 172 -1018
rect 146 -1023 150 -1019
rect 168 -1023 172 -1019
rect 178 -1023 182 -1018
rect 197 -1018 211 -1014
rect 219 -1018 255 -1015
rect 157 -1046 161 -1043
rect 190 -1046 194 -1043
rect 197 -1046 200 -1018
rect 219 -1019 245 -1018
rect 219 -1023 223 -1019
rect 241 -1023 245 -1019
rect 251 -1023 255 -1018
rect 270 -1018 292 -1014
rect 157 -1050 181 -1046
rect 190 -1050 200 -1046
rect 230 -1046 234 -1043
rect 263 -1046 267 -1043
rect 270 -1046 273 -1018
rect 376 -1019 379 -991
rect 420 -1006 426 -1002
rect 412 -1019 415 -1016
rect 420 -1019 423 -1006
rect 438 -1006 444 -1002
rect 578 -988 582 -983
rect 287 -1024 320 -1021
rect 287 -1025 294 -1024
rect 230 -1050 254 -1046
rect 263 -1050 273 -1046
rect 290 -1028 294 -1025
rect 316 -1028 320 -1024
rect 412 -1022 423 -1019
rect 137 -1055 147 -1051
rect 137 -1084 140 -1055
rect 160 -1057 161 -1053
rect 168 -1058 172 -1050
rect 190 -1058 194 -1050
rect 213 -1055 220 -1051
rect 146 -1074 150 -1068
rect 178 -1074 182 -1068
rect 146 -1077 182 -1074
rect 163 -1081 170 -1077
rect 213 -1084 216 -1055
rect 233 -1057 234 -1053
rect 241 -1058 245 -1050
rect 263 -1058 267 -1050
rect 307 -1051 311 -1048
rect 324 -1051 328 -1048
rect 299 -1055 317 -1051
rect 324 -1054 335 -1051
rect 299 -1060 303 -1055
rect 324 -1060 328 -1054
rect 219 -1074 223 -1068
rect 251 -1074 255 -1068
rect 219 -1077 255 -1074
rect 290 -1074 294 -1070
rect 308 -1074 312 -1070
rect 316 -1074 320 -1070
rect 290 -1077 320 -1074
rect 236 -1081 243 -1077
rect 303 -1080 306 -1077
rect 137 -1087 216 -1084
rect 137 -1143 141 -1087
rect 331 -1106 335 -1054
rect 144 -1110 180 -1107
rect 144 -1111 170 -1110
rect 144 -1115 148 -1111
rect 166 -1115 170 -1111
rect 176 -1115 180 -1110
rect 195 -1110 211 -1106
rect 228 -1110 335 -1106
rect 376 -1095 379 -1024
rect 420 -1031 423 -1022
rect 441 -1019 444 -1006
rect 495 -1008 499 -1005
rect 450 -1012 488 -1008
rect 495 -1012 505 -1008
rect 450 -1019 453 -1012
rect 495 -1017 499 -1012
rect 441 -1022 453 -1019
rect 420 -1035 426 -1031
rect 441 -1031 444 -1022
rect 438 -1035 444 -1031
rect 420 -1045 427 -1041
rect 396 -1067 404 -1064
rect 399 -1072 403 -1067
rect 376 -1099 400 -1095
rect 407 -1096 411 -1092
rect 420 -1074 424 -1045
rect 450 -1054 453 -1022
rect 502 -1022 505 -1012
rect 511 -1013 517 -1009
rect 511 -1022 514 -1013
rect 529 -1013 535 -1009
rect 586 -1011 590 -1008
rect 502 -1025 514 -1022
rect 457 -1034 463 -1030
rect 457 -1054 460 -1034
rect 475 -1034 481 -1030
rect 450 -1057 460 -1054
rect 457 -1059 460 -1057
rect 457 -1063 463 -1059
rect 478 -1057 481 -1034
rect 487 -1033 491 -1027
rect 487 -1036 499 -1033
rect 495 -1042 499 -1036
rect 487 -1057 491 -1052
rect 502 -1056 505 -1025
rect 511 -1038 514 -1025
rect 532 -1029 535 -1013
rect 541 -1015 579 -1011
rect 586 -1015 596 -1011
rect 541 -1029 544 -1015
rect 586 -1020 590 -1015
rect 511 -1042 517 -1038
rect 532 -1033 544 -1029
rect 532 -1038 535 -1033
rect 529 -1042 535 -1038
rect 501 -1057 505 -1056
rect 478 -1059 491 -1057
rect 475 -1061 491 -1059
rect 498 -1061 505 -1057
rect 511 -1057 518 -1053
rect 541 -1057 544 -1033
rect 593 -1021 596 -1015
rect 593 -1024 607 -1021
rect 578 -1036 582 -1030
rect 578 -1039 590 -1036
rect 548 -1055 554 -1051
rect 548 -1057 551 -1055
rect 475 -1063 481 -1061
rect 487 -1064 491 -1061
rect 420 -1078 464 -1074
rect 420 -1096 424 -1078
rect 495 -1089 499 -1084
rect 494 -1092 502 -1089
rect 511 -1090 515 -1057
rect 541 -1060 551 -1057
rect 548 -1080 551 -1060
rect 586 -1045 590 -1039
rect 566 -1055 572 -1051
rect 569 -1060 572 -1055
rect 578 -1060 582 -1055
rect 593 -1059 596 -1024
rect 592 -1060 596 -1059
rect 569 -1064 582 -1060
rect 589 -1064 596 -1060
rect 548 -1084 554 -1080
rect 569 -1080 572 -1064
rect 566 -1084 572 -1080
rect 578 -1067 582 -1064
rect 511 -1094 555 -1090
rect 586 -1092 590 -1087
rect 511 -1096 516 -1094
rect 585 -1095 593 -1092
rect 407 -1097 412 -1096
rect 420 -1097 516 -1096
rect 155 -1138 159 -1135
rect 188 -1138 192 -1135
rect 195 -1138 198 -1110
rect 206 -1116 239 -1113
rect 206 -1117 213 -1116
rect 155 -1142 179 -1138
rect 188 -1142 198 -1138
rect 209 -1120 213 -1117
rect 235 -1120 239 -1116
rect 251 -1117 261 -1113
rect 278 -1117 315 -1113
rect 137 -1147 145 -1143
rect 158 -1149 159 -1145
rect 166 -1150 170 -1142
rect 188 -1150 192 -1142
rect 226 -1143 230 -1140
rect 243 -1143 247 -1140
rect 251 -1143 254 -1117
rect 218 -1147 236 -1143
rect 243 -1146 254 -1143
rect 259 -1123 289 -1120
rect 259 -1127 263 -1123
rect 285 -1127 289 -1123
rect 218 -1152 222 -1147
rect 243 -1152 247 -1146
rect 276 -1150 280 -1147
rect 144 -1166 148 -1160
rect 176 -1166 180 -1160
rect 144 -1169 180 -1166
rect 209 -1166 213 -1162
rect 227 -1166 231 -1162
rect 268 -1154 286 -1150
rect 268 -1159 272 -1154
rect 293 -1159 297 -1147
rect 235 -1166 239 -1162
rect 209 -1169 239 -1166
rect 161 -1173 168 -1169
rect 222 -1172 225 -1169
rect 259 -1173 263 -1169
rect 277 -1173 281 -1169
rect 285 -1173 289 -1169
rect 259 -1176 289 -1173
rect 272 -1179 275 -1176
rect 312 -1194 315 -1117
rect 85 -1197 315 -1194
rect 376 -1215 379 -1099
rect 407 -1100 516 -1097
rect 407 -1104 411 -1100
rect 399 -1119 403 -1114
rect -282 -1219 379 -1215
<< m2contact >>
rect -292 61 -287 66
rect -142 73 -136 79
rect -244 61 -239 66
rect -278 52 -273 57
rect -195 52 -190 57
rect -104 36 -99 41
rect -292 -81 -287 -76
rect -244 -81 -239 -76
rect -142 -68 -136 -62
rect -278 -89 -273 -84
rect -195 -89 -190 -84
rect 123 40 128 45
rect 123 -6 128 -1
rect -23 -19 -18 -14
rect -104 -105 -99 -100
rect -23 -36 -18 -31
rect 289 6 294 11
rect 362 16 367 21
rect 318 6 323 11
rect 410 16 415 21
rect 512 29 518 35
rect 376 8 381 13
rect 459 8 464 13
rect 550 -8 555 -3
rect 35 -120 40 -115
rect 35 -147 40 -142
rect 202 -166 207 -161
rect -293 -226 -288 -221
rect -245 -226 -240 -221
rect -143 -214 -137 -208
rect -279 -235 -274 -230
rect -196 -235 -191 -230
rect -105 -251 -100 -246
rect -293 -368 -288 -363
rect -245 -368 -240 -363
rect -143 -355 -137 -349
rect -279 -376 -274 -371
rect -196 -376 -191 -371
rect -24 -268 -19 -263
rect -105 -392 -100 -387
rect -24 -285 -19 -280
rect 34 -369 39 -364
rect 34 -396 39 -391
rect 256 -243 261 -238
rect 298 -166 303 -161
rect 410 -244 415 -239
rect 512 -231 518 -225
rect 376 -252 381 -247
rect 459 -252 464 -247
rect 550 -268 555 -263
rect 149 -347 154 -342
rect 191 -385 196 -380
rect 149 -393 154 -388
rect 255 -390 260 -385
rect 255 -443 260 -438
rect -294 -510 -289 -505
rect -246 -510 -241 -505
rect -144 -498 -138 -492
rect -280 -519 -275 -514
rect -197 -519 -192 -514
rect -106 -535 -101 -530
rect -294 -652 -289 -647
rect -246 -652 -241 -647
rect -144 -639 -138 -633
rect -280 -660 -275 -655
rect -197 -660 -192 -655
rect -18 -553 -13 -548
rect -106 -676 -101 -671
rect -18 -570 -13 -565
rect 40 -654 45 -649
rect 40 -681 45 -676
rect -294 -799 -289 -794
rect -246 -799 -241 -794
rect -144 -787 -138 -781
rect -280 -808 -275 -803
rect -197 -808 -192 -803
rect 262 -528 267 -523
rect 410 -528 415 -523
rect 512 -515 518 -509
rect 376 -536 381 -531
rect 459 -536 464 -531
rect 550 -552 555 -547
rect 155 -632 160 -627
rect 197 -670 203 -664
rect 270 -670 275 -665
rect 155 -678 160 -673
rect 228 -678 233 -673
rect 284 -756 289 -751
rect -106 -824 -101 -819
rect 284 -809 289 -804
rect -294 -941 -289 -936
rect -246 -941 -241 -936
rect -144 -928 -138 -922
rect -280 -949 -275 -944
rect -197 -949 -192 -944
rect -18 -915 -13 -910
rect -18 -933 -13 -928
rect -106 -965 -101 -960
rect -29 -984 -24 -979
rect -18 -950 -13 -945
rect 47 -915 52 -910
rect 142 -908 147 -903
rect 47 -984 52 -979
rect 40 -1034 45 -1029
rect 40 -1061 45 -1056
rect 204 -908 209 -903
rect 262 -908 267 -903
rect 291 -908 296 -903
rect 328 -908 333 -903
rect 410 -797 415 -792
rect 512 -784 518 -778
rect 376 -805 381 -800
rect 459 -805 464 -800
rect 550 -821 555 -816
rect 155 -1012 160 -1007
rect 410 -1016 415 -1011
rect 512 -1003 518 -997
rect 376 -1024 381 -1019
rect 155 -1058 160 -1053
rect 228 -1058 233 -1053
rect 459 -1024 464 -1019
rect 550 -1040 555 -1035
rect 153 -1150 158 -1145
rect 297 -1155 302 -1150
<< metal2 >>
rect -150 83 -100 86
rect -150 78 -147 83
rect -202 75 -142 78
rect -287 62 -244 65
rect -202 56 -199 75
rect -273 53 -195 56
rect -103 41 -100 83
rect 123 -1 128 40
rect 504 39 554 42
rect 504 34 507 39
rect 452 31 512 34
rect 367 17 410 20
rect 294 7 318 10
rect 452 12 455 31
rect 381 9 459 12
rect 551 -3 554 39
rect -23 -31 -18 -19
rect -150 -58 -100 -55
rect -150 -63 -147 -58
rect -202 -66 -142 -63
rect -287 -80 -244 -77
rect -202 -85 -199 -66
rect -273 -88 -195 -85
rect -103 -100 -100 -58
rect 35 -142 40 -120
rect 207 -166 298 -161
rect -151 -204 -101 -201
rect -151 -209 -148 -204
rect -203 -212 -143 -209
rect -288 -225 -245 -222
rect -203 -231 -200 -212
rect -274 -234 -196 -231
rect -104 -246 -101 -204
rect 504 -221 554 -218
rect 504 -226 507 -221
rect 452 -229 512 -226
rect 369 -239 372 -238
rect 261 -240 372 -239
rect 261 -242 410 -240
rect 369 -243 410 -242
rect 452 -248 455 -229
rect 381 -251 459 -248
rect 551 -263 554 -221
rect -24 -280 -19 -268
rect -151 -345 -101 -342
rect -151 -350 -148 -345
rect -203 -353 -143 -350
rect -288 -367 -245 -364
rect -203 -372 -200 -353
rect -274 -375 -196 -372
rect -104 -387 -101 -345
rect 34 -391 39 -369
rect 149 -388 154 -347
rect 191 -453 196 -385
rect 255 -438 260 -390
rect 191 -456 233 -453
rect -152 -488 -102 -485
rect -152 -493 -149 -488
rect -204 -496 -144 -493
rect -289 -509 -246 -506
rect -204 -515 -201 -496
rect -275 -518 -197 -515
rect -105 -530 -102 -488
rect -18 -565 -13 -553
rect -152 -629 -102 -626
rect -152 -634 -149 -629
rect -204 -637 -144 -634
rect -289 -651 -246 -648
rect -204 -656 -201 -637
rect -275 -659 -197 -656
rect -105 -671 -102 -629
rect 40 -676 45 -654
rect 155 -673 160 -632
rect -152 -777 -102 -774
rect -152 -782 -149 -777
rect -204 -785 -144 -782
rect -289 -798 -246 -795
rect -204 -804 -201 -785
rect -275 -807 -197 -804
rect -105 -819 -102 -777
rect 198 -838 201 -670
rect 228 -673 233 -456
rect 504 -505 554 -502
rect 504 -510 507 -505
rect 452 -513 512 -510
rect 267 -527 410 -524
rect 452 -532 455 -513
rect 381 -535 459 -532
rect 551 -547 554 -505
rect 198 -842 233 -838
rect 147 -907 155 -904
rect 202 -907 204 -904
rect -13 -914 47 -911
rect -152 -918 -102 -915
rect -152 -923 -149 -918
rect -204 -926 -144 -923
rect -289 -940 -246 -937
rect -204 -945 -201 -926
rect -275 -948 -197 -945
rect -105 -960 -102 -918
rect -18 -945 -13 -933
rect -24 -983 47 -980
rect 40 -1056 45 -1034
rect 155 -1053 160 -1012
rect 228 -1053 233 -842
rect 271 -894 274 -670
rect 284 -804 289 -756
rect 504 -774 554 -771
rect 504 -779 507 -774
rect 452 -782 512 -779
rect 329 -796 410 -793
rect 271 -897 303 -894
rect 267 -907 291 -904
rect 300 -931 303 -897
rect 329 -903 332 -796
rect 452 -801 455 -782
rect 381 -804 459 -801
rect 551 -816 554 -774
rect 250 -934 303 -931
rect 250 -1101 253 -934
rect 504 -993 554 -990
rect 504 -998 507 -993
rect 452 -1001 512 -998
rect 153 -1104 253 -1101
rect 348 -1015 410 -1012
rect 153 -1145 158 -1104
rect 348 -1151 351 -1015
rect 452 -1020 455 -1001
rect 381 -1023 459 -1020
rect 551 -1035 554 -993
rect 302 -1154 351 -1151
use dff  dff_0
timestamp 1618572623
transform 1 0 -129 0 1 -49
box -131 6 76 148
use xor  xor_0
timestamp 1618484725
transform 1 0 0 0 1 -22
box -11 -51 105 80
use and  and_1
timestamp 1618590203
transform 1 0 111 0 1 -25
box 1 0 54 62
use xor  xor_1
timestamp 1618484725
transform 1 0 189 0 1 -15
box -11 -51 105 80
use and  and_0
timestamp 1618590203
transform 1 0 22 0 1 -139
box 1 0 54 62
use or  or_0
timestamp 1618732609
transform 1 0 118 0 1 -112
box -27 -27 14 35
<< labels >>
rlabel metal1 -39 35 -39 35 3 a1
rlabel metal1 -38 26 -38 26 3 b1
rlabel metal1 46 2 46 2 1 a1
rlabel metal1 46 -67 46 -67 1 b1
rlabel metal1 110 1 110 1 1 p1
rlabel metal1 166 4 166 4 1 i1
rlabel metal1 77 -110 77 -110 1 g1
rlabel metal1 235 9 235 9 1 p1
rlabel metal1 325 9 325 9 7 sum1
rlabel metal1 125 46 125 46 1 c0
rlabel metal1 312 75 312 75 5 c0
rlabel metal1 -40 -213 -40 -213 3 a2
rlabel metal1 -37 -222 -37 -222 1 b2
rlabel metal1 42 -194 42 -194 1 vdd
rlabel metal1 45 -262 45 -262 1 vdd
rlabel metal1 34 -250 34 -250 1 gnd
rlabel metal1 -8 -261 -8 -261 1 gnd
rlabel metal1 70 -274 70 -274 1 gnd
rlabel metal1 33 -318 33 -318 1 gnd
rlabel metal1 25 -385 25 -385 1 gnd
rlabel metal1 37 -328 37 -328 1 vdd
rlabel metal1 45 -247 45 -247 1 a2
rlabel metal1 45 -316 45 -316 1 b2
rlabel metal1 99 -248 99 -248 1 p2
rlabel metal1 74 -359 74 -359 1 g2
rlabel metal1 41 61 41 61 1 vdd
rlabel metal1 51 -10 51 -10 1 vdd
rlabel metal1 46 -76 46 -76 1 vdd
rlabel metal1 113 36 113 36 1 vdd
rlabel metal1 231 66 231 66 1 vdd
rlabel metal1 239 -2 239 -2 1 vdd
rlabel metal1 34 -7 34 -7 1 gnd
rlabel metal1 72 -28 72 -28 1 gnd
rlabel metal1 -12 -10 -12 -10 1 gnd
rlabel metal1 54 -140 54 -140 1 gnd
rlabel metal1 106 -140 106 -140 1 gnd
rlabel metal1 136 -28 136 -28 1 gnd
rlabel metal1 180 -1 180 -1 1 gnd
rlabel metal1 90 -85 90 -85 1 vdd
rlabel metal1 226 3 226 3 1 gnd
rlabel metal1 260 -21 260 -21 1 gnd
rlabel metal1 215 -64 215 -64 1 gnd
rlabel metal1 205 -186 205 -186 1 vdd
rlabel metal1 202 -253 202 -253 1 vdd
rlabel metal1 189 -313 189 -313 1 gnd
rlabel metal1 149 -253 149 -253 1 gnd
rlabel metal1 191 -246 191 -246 1 gnd
rlabel metal1 229 -268 229 -268 1 gnd
rlabel metal1 202 -240 202 -240 1 p2
rlabel metal1 142 -351 142 -351 1 vdd
rlabel metal1 160 -414 160 -414 1 gnd
rlabel metal1 228 -414 228 -414 1 gnd
rlabel metal1 236 -358 236 -358 1 vdd
rlabel metal1 253 -387 253 -387 1 c2
rlabel metal1 48 -479 48 -479 1 vdd
rlabel metal1 51 -547 51 -547 1 vdd
rlabel metal1 40 -535 40 -535 1 gnd
rlabel metal1 -2 -546 -2 -546 1 gnd
rlabel metal1 76 -559 76 -559 1 gnd
rlabel metal1 39 -603 39 -603 1 gnd
rlabel metal1 31 -670 31 -670 1 gnd
rlabel metal1 43 -613 43 -613 1 vdd
rlabel metal1 211 -471 211 -471 1 vdd
rlabel metal1 208 -538 208 -538 1 vdd
rlabel metal1 195 -598 195 -598 1 gnd
rlabel metal1 155 -538 155 -538 1 gnd
rlabel metal1 197 -531 197 -531 1 gnd
rlabel metal1 235 -553 235 -553 1 gnd
rlabel metal1 148 -636 148 -636 1 vdd
rlabel metal1 166 -699 166 -699 1 gnd
rlabel metal1 -30 -499 -30 -499 1 a3
rlabel metal1 -32 -508 -32 -508 1 b3
rlabel metal1 51 -532 51 -532 1 a3
rlabel metal1 51 -602 51 -602 1 b3
rlabel metal1 113 -532 113 -532 1 p3
rlabel metal1 136 -114 136 -114 1 c1
rlabel metal1 239 -699 239 -699 1 gnd
rlabel metal1 221 -636 221 -636 1 vdd
rlabel metal1 304 -699 304 -699 1 gnd
rlabel metal1 312 -643 312 -643 1 vdd
rlabel metal1 257 -780 257 -780 1 gnd
rlabel metal1 265 -724 265 -724 1 vdd
rlabel metal1 282 -754 282 -754 1 c3
rlabel metal1 208 -524 208 -524 1 p3
rlabel metal1 48 -859 48 -859 1 vdd
rlabel metal1 51 -927 51 -927 1 vdd
rlabel metal1 40 -915 40 -915 1 gnd
rlabel metal1 -2 -926 -2 -926 1 gnd
rlabel metal1 76 -939 76 -939 1 gnd
rlabel metal1 39 -983 39 -983 1 gnd
rlabel metal1 31 -1050 31 -1050 1 gnd
rlabel metal1 43 -993 43 -993 1 vdd
rlabel metal1 211 -851 211 -851 1 vdd
rlabel metal1 208 -918 208 -918 1 vdd
rlabel metal1 195 -978 195 -978 1 gnd
rlabel metal1 155 -918 155 -918 1 gnd
rlabel metal1 197 -911 197 -911 1 gnd
rlabel metal1 235 -933 235 -933 1 gnd
rlabel metal1 148 -1016 148 -1016 1 vdd
rlabel metal1 166 -1079 166 -1079 1 gnd
rlabel metal1 239 -1079 239 -1079 1 gnd
rlabel metal1 221 -1016 221 -1016 1 vdd
rlabel metal1 -33 -878 -33 -878 1 a4
rlabel metal1 -33 -887 -33 -887 1 b4
rlabel metal1 116 -913 116 -913 1 p4
rlabel metal1 82 -1025 82 -1025 1 g4
rlabel metal1 81 -645 81 -645 1 g3
rlabel metal1 146 -1108 146 -1108 1 vdd
rlabel metal1 164 -1171 164 -1171 1 gnd
rlabel metal1 305 -1079 305 -1079 1 gnd
rlabel metal1 313 -1023 313 -1023 1 vdd
rlabel metal1 224 -1171 224 -1171 1 gnd
rlabel metal1 232 -1115 232 -1115 1 vdd
rlabel metal1 274 -1178 274 -1178 1 gnd
rlabel metal1 282 -1122 282 -1122 1 vdd
rlabel metal2 203 -906 203 -906 1 p4
rlabel m2contact -138 -67 -138 -67 1 clk
rlabel m2contact -101 -103 -101 -103 3 clk
rlabel metal1 -66 -158 -66 -158 1 vdd
rlabel metal1 -67 -103 -67 -103 1 gnd
rlabel metal1 -76 -46 -76 -46 5 vdd
rlabel m2contact -191 -88 -191 -88 1 clk
rlabel metal1 -228 -54 -228 -54 1 clk
rlabel metal1 -167 -43 -167 -43 5 vdd
rlabel metal1 -158 -100 -158 -100 1 gnd
rlabel metal1 -157 -155 -157 -155 1 vdd
rlabel metal1 -253 -182 -253 -182 1 gnd
rlabel metal1 -253 -131 -253 -131 1 vdd
rlabel metal1 -257 -162 -257 -162 3 clk
rlabel metal1 -295 -78 -295 -78 3 bin1
rlabel metal1 -294 63 -294 63 3 ain1
rlabel metal1 -277 98 -277 98 5 clk
rlabel m2contact -139 -354 -139 -354 1 clk
rlabel m2contact -102 -390 -102 -390 3 clk
rlabel metal1 -67 -445 -67 -445 1 vdd
rlabel metal1 -68 -390 -68 -390 1 gnd
rlabel metal1 -77 -333 -77 -333 5 vdd
rlabel m2contact -192 -375 -192 -375 1 clk
rlabel metal1 -229 -341 -229 -341 1 clk
rlabel metal1 -168 -330 -168 -330 5 vdd
rlabel metal1 -159 -387 -159 -387 1 gnd
rlabel metal1 -158 -442 -158 -442 1 vdd
rlabel metal1 -254 -469 -254 -469 1 gnd
rlabel metal1 -254 -418 -254 -418 1 vdd
rlabel metal1 -258 -449 -258 -449 3 clk
rlabel metal1 -278 -189 -278 -189 5 clk
rlabel metal1 -258 -308 -258 -308 3 clk
rlabel metal1 -254 -277 -254 -277 1 vdd
rlabel metal1 -254 -328 -254 -328 1 gnd
rlabel metal1 -158 -301 -158 -301 1 vdd
rlabel metal1 -159 -246 -159 -246 1 gnd
rlabel metal1 -168 -189 -168 -189 5 vdd
rlabel metal1 -229 -200 -229 -200 1 clk
rlabel m2contact -192 -234 -192 -234 1 clk
rlabel metal1 -77 -192 -77 -192 5 vdd
rlabel metal1 -68 -249 -68 -249 1 gnd
rlabel metal1 -67 -304 -67 -304 1 vdd
rlabel m2contact -102 -249 -102 -249 3 clk
rlabel m2contact -139 -213 -139 -213 1 clk
rlabel metal1 -296 -366 -296 -366 3 bin2
rlabel metal1 -297 -650 -297 -650 3 bin3
rlabel m2contact -140 -638 -140 -638 1 clk
rlabel m2contact -103 -674 -103 -674 3 clk
rlabel metal1 -68 -729 -68 -729 1 vdd
rlabel metal1 -69 -674 -69 -674 1 gnd
rlabel metal1 -78 -617 -78 -617 5 vdd
rlabel m2contact -193 -659 -193 -659 1 clk
rlabel metal1 -230 -625 -230 -625 1 clk
rlabel metal1 -169 -614 -169 -614 5 vdd
rlabel metal1 -160 -671 -160 -671 1 gnd
rlabel metal1 -159 -726 -159 -726 1 vdd
rlabel metal1 -255 -753 -255 -753 1 gnd
rlabel metal1 -255 -702 -255 -702 1 vdd
rlabel metal1 -259 -733 -259 -733 3 clk
rlabel metal1 -279 -473 -279 -473 5 clk
rlabel metal1 -259 -592 -259 -592 3 clk
rlabel metal1 -255 -561 -255 -561 1 vdd
rlabel metal1 -255 -612 -255 -612 1 gnd
rlabel metal1 -159 -585 -159 -585 1 vdd
rlabel metal1 -160 -530 -160 -530 1 gnd
rlabel metal1 -169 -473 -169 -473 5 vdd
rlabel metal1 -230 -484 -230 -484 1 clk
rlabel m2contact -193 -518 -193 -518 1 clk
rlabel metal1 -78 -476 -78 -476 5 vdd
rlabel metal1 -69 -533 -69 -533 1 gnd
rlabel metal1 -68 -588 -68 -588 1 vdd
rlabel m2contact -103 -533 -103 -533 3 clk
rlabel m2contact -140 -497 -140 -497 1 clk
rlabel m2contact -140 -927 -140 -927 1 clk
rlabel m2contact -103 -963 -103 -963 3 clk
rlabel metal1 -68 -1018 -68 -1018 1 vdd
rlabel metal1 -69 -963 -69 -963 1 gnd
rlabel metal1 -78 -906 -78 -906 5 vdd
rlabel m2contact -193 -948 -193 -948 1 clk
rlabel metal1 -230 -914 -230 -914 1 clk
rlabel metal1 -169 -903 -169 -903 5 vdd
rlabel metal1 -160 -960 -160 -960 1 gnd
rlabel metal1 -159 -1015 -159 -1015 1 vdd
rlabel metal1 -255 -1042 -255 -1042 1 gnd
rlabel metal1 -255 -991 -255 -991 1 vdd
rlabel metal1 -259 -1022 -259 -1022 3 clk
rlabel metal1 -279 -762 -279 -762 5 clk
rlabel metal1 -259 -881 -259 -881 3 clk
rlabel metal1 -255 -850 -255 -850 1 vdd
rlabel metal1 -255 -901 -255 -901 1 gnd
rlabel metal1 -159 -874 -159 -874 1 vdd
rlabel metal1 -160 -819 -160 -819 1 gnd
rlabel metal1 -169 -762 -169 -762 5 vdd
rlabel metal1 -230 -773 -230 -773 1 clk
rlabel m2contact -193 -807 -193 -807 1 clk
rlabel metal1 -78 -765 -78 -765 5 vdd
rlabel metal1 -69 -822 -69 -822 1 gnd
rlabel metal1 -68 -877 -68 -877 1 vdd
rlabel m2contact -103 -822 -103 -822 3 clk
rlabel m2contact -140 -786 -140 -786 1 clk
rlabel metal1 -296 -938 -296 -938 3 bin4
rlabel metal1 -297 -508 -297 -508 3 ain3
rlabel metal1 -296 -797 -296 -797 3 ain4
rlabel metal1 -295 -224 -295 -224 3 ain2
rlabel metal1 -165 100 -165 100 5 vdd
rlabel metal1 -74 97 -74 97 5 vdd
rlabel metal1 -253 13 -253 13 1 vdd
rlabel metal1 -151 -15 -151 -15 1 vdd
rlabel metal1 -60 -17 -60 -17 1 vdd
rlabel metal1 -253 -44 -253 -44 1 gnd
rlabel metal1 -168 41 -168 41 1 gnd
rlabel metal1 -77 38 -77 38 1 gnd
rlabel metal1 397 -65 397 -65 3 clk
rlabel metal1 401 -34 401 -34 1 vdd
rlabel metal1 401 -85 401 -85 1 gnd
rlabel metal1 497 -58 497 -58 1 vdd
rlabel metal1 496 -3 496 -3 1 gnd
rlabel metal1 487 54 487 54 5 vdd
rlabel metal1 426 43 426 43 1 clk
rlabel m2contact 463 9 463 9 1 clk
rlabel metal1 578 51 578 51 5 vdd
rlabel metal1 587 -6 587 -6 1 gnd
rlabel metal1 588 -61 588 -61 1 vdd
rlabel m2contact 553 -6 553 -6 3 clk
rlabel m2contact 516 30 516 30 1 clk
rlabel metal1 601 10 601 10 1 sum1out
rlabel metal1 254 -241 254 -241 1 sum2
rlabel m2contact 516 -230 516 -230 1 clk
rlabel m2contact 553 -266 553 -266 3 clk
rlabel metal1 588 -321 588 -321 1 vdd
rlabel metal1 587 -266 587 -266 1 gnd
rlabel metal1 578 -209 578 -209 5 vdd
rlabel m2contact 463 -251 463 -251 1 clk
rlabel metal1 426 -217 426 -217 1 clk
rlabel metal1 487 -206 487 -206 5 vdd
rlabel metal1 496 -263 496 -263 1 gnd
rlabel metal1 497 -318 497 -318 1 vdd
rlabel metal1 401 -345 401 -345 1 gnd
rlabel metal1 401 -294 401 -294 1 vdd
rlabel metal1 397 -325 397 -325 3 clk
rlabel metal1 601 -250 601 -250 1 sum2out
rlabel metal1 259 -526 259 -526 1 sum3
rlabel metal1 397 -609 397 -609 3 clk
rlabel metal1 401 -578 401 -578 1 vdd
rlabel metal1 401 -629 401 -629 1 gnd
rlabel metal1 497 -602 497 -602 1 vdd
rlabel metal1 496 -547 496 -547 1 gnd
rlabel metal1 487 -490 487 -490 5 vdd
rlabel metal1 426 -501 426 -501 1 clk
rlabel m2contact 463 -535 463 -535 1 clk
rlabel metal1 578 -493 578 -493 5 vdd
rlabel metal1 587 -550 587 -550 1 gnd
rlabel metal1 588 -605 588 -605 1 vdd
rlabel m2contact 553 -550 553 -550 3 clk
rlabel m2contact 516 -514 516 -514 1 clk
rlabel metal1 604 -534 604 -534 7 sum3out
rlabel metal1 397 -878 397 -878 3 clk
rlabel metal1 401 -847 401 -847 1 vdd
rlabel metal1 401 -898 401 -898 1 gnd
rlabel metal1 497 -871 497 -871 1 vdd
rlabel metal1 496 -816 496 -816 1 gnd
rlabel metal1 487 -759 487 -759 5 vdd
rlabel metal1 426 -770 426 -770 1 clk
rlabel m2contact 463 -804 463 -804 1 clk
rlabel metal1 578 -762 578 -762 5 vdd
rlabel metal1 587 -819 587 -819 1 gnd
rlabel metal1 588 -874 588 -874 1 vdd
rlabel m2contact 553 -819 553 -819 3 clk
rlabel m2contact 516 -783 516 -783 1 clk
rlabel metal1 260 -905 260 -905 1 sum4
rlabel metal1 397 -1097 397 -1097 3 clk
rlabel metal1 401 -1066 401 -1066 1 vdd
rlabel metal1 401 -1117 401 -1117 1 gnd
rlabel metal1 497 -1090 497 -1090 1 vdd
rlabel metal1 496 -1035 496 -1035 1 gnd
rlabel metal1 487 -978 487 -978 5 vdd
rlabel metal1 426 -989 426 -989 1 clk
rlabel m2contact 463 -1023 463 -1023 1 clk
rlabel metal1 578 -981 578 -981 5 vdd
rlabel metal1 587 -1038 587 -1038 1 gnd
rlabel metal1 588 -1093 588 -1093 1 vdd
rlabel m2contact 553 -1038 553 -1038 3 clk
rlabel m2contact 516 -1002 516 -1002 1 clk
rlabel metal1 295 -1152 295 -1152 1 cout
rlabel metal1 603 -802 603 -802 7 sum4out
rlabel metal1 604 -1022 604 -1022 7 cout_out
<< end >>
