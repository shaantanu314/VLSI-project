magic
tech scmos
timestamp 1618406033
<< ntransistor >>
rect -4 -25 -2 -15
rect 10 -25 12 -15
<< ptransistor >>
rect -4 0 -2 20
rect 10 0 12 20
<< ndiffusion >>
rect -5 -25 -4 -15
rect -2 -25 10 -15
rect 12 -25 13 -15
<< pdiffusion >>
rect -5 0 -4 20
rect -2 0 2 20
rect 6 0 10 20
rect 12 0 13 20
<< ndcontact >>
rect -9 -25 -5 -15
rect 13 -25 17 -15
<< pdcontact >>
rect -9 0 -5 20
rect 2 0 6 20
rect 13 0 17 20
<< polysilicon >>
rect -4 20 -2 23
rect 10 20 12 23
rect -4 -15 -2 0
rect 10 -15 12 0
rect -4 -30 -2 -25
rect 10 -30 12 -25
<< metal1 >>
rect -9 24 17 28
rect -9 20 -5 24
rect 13 20 17 24
rect 2 -3 6 0
rect 2 -7 18 -3
rect 13 -15 17 -7
rect -9 -30 -5 -25
rect -11 -34 -5 -30
<< labels >>
rlabel metal1 4 27 4 27 5 vdd
rlabel metal1 16 -5 16 -5 7 out
rlabel metal1 -8 -32 -8 -32 2 gnd
<< end >>
