magic
tech scmos
timestamp 1613754354
<< nwell >>
rect 0 0 24 37
<< ntransistor >>
rect 11 -18 13 -8
<< ptransistor >>
rect 11 6 13 31
<< ndiffusion >>
rect 10 -18 11 -8
rect 13 -18 14 -8
<< pdiffusion >>
rect 10 6 11 31
rect 13 6 14 31
<< ndcontact >>
rect 6 -18 10 -8
rect 14 -18 18 -8
<< pdcontact >>
rect 6 6 10 31
rect 14 6 18 31
<< polysilicon >>
rect 11 31 13 34
rect 11 -8 13 6
rect 11 -21 13 -18
<< polycontact >>
rect 7 -5 11 -1
<< metal1 >>
rect 0 36 24 40
rect 6 31 10 36
rect 14 -1 18 6
rect -3 -5 7 -1
rect 14 -5 27 -1
rect 14 -8 18 -5
rect 6 -24 10 -18
rect 0 -28 24 -24
<< labels >>
flabel metal1 -3 -5 7 -1 7 FreeSans 23 0 0 0 in
flabel metal1 14 -5 27 -1 3 FreeSans 23 0 8 0 out
flabel space -2 5 25 32 3 FreeSans 23 0 52 0 pmos
flabel space 0 -19 22 -7 3 FreeSans 23 0 56 0 nmos
rlabel metal1 0 -28 24 -24 1 gnd
rlabel metal1 0 36 24 40 5 vdd
rlabel space 6 -18 18 -8 1 gnd
<< end >>
