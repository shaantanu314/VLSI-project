magic
tech scmos
timestamp 1619416395
<< ntransistor >>
rect -3 -253 -1 -243
rect 11 -253 13 -243
rect 36 -244 38 -234
rect 50 -244 52 -234
rect 154 -246 156 -236
rect 168 -246 170 -236
rect 193 -237 195 -227
rect 207 -237 209 -227
rect 76 -267 78 -257
rect 90 -267 92 -257
rect 233 -260 235 -250
rect 247 -260 249 -250
rect 36 -313 38 -303
rect 50 -313 52 -303
rect 193 -306 195 -296
rect 207 -306 209 -296
rect 29 -379 31 -369
rect 43 -379 45 -369
rect 63 -379 65 -369
rect 145 -403 147 -393
rect 159 -403 161 -393
rect 179 -403 181 -393
rect 219 -405 221 -395
rect 227 -405 229 -395
rect 244 -405 246 -395
rect 3 -538 5 -528
rect 17 -538 19 -528
rect 42 -529 44 -519
rect 56 -529 58 -519
rect 160 -531 162 -521
rect 174 -531 176 -521
rect 199 -522 201 -512
rect 213 -522 215 -512
rect 82 -552 84 -542
rect 96 -552 98 -542
rect 239 -545 241 -535
rect 253 -545 255 -535
rect 42 -598 44 -588
rect 56 -598 58 -588
rect 199 -591 201 -581
rect 213 -591 215 -581
rect 35 -664 37 -654
rect 49 -664 51 -654
rect 69 -664 71 -654
rect 151 -688 153 -678
rect 165 -688 167 -678
rect 185 -688 187 -678
rect 224 -688 226 -678
rect 238 -688 240 -678
rect 258 -688 260 -678
rect 295 -690 297 -680
rect 303 -690 305 -680
rect 320 -690 322 -680
rect 248 -771 250 -761
rect 256 -771 258 -761
rect 273 -771 275 -761
rect 3 -918 5 -908
rect 17 -918 19 -908
rect 42 -909 44 -899
rect 56 -909 58 -899
rect 160 -911 162 -901
rect 174 -911 176 -901
rect 199 -902 201 -892
rect 213 -902 215 -892
rect 82 -932 84 -922
rect 96 -932 98 -922
rect 239 -925 241 -915
rect 253 -925 255 -915
rect 42 -978 44 -968
rect 56 -978 58 -968
rect 199 -971 201 -961
rect 213 -971 215 -961
rect 35 -1044 37 -1034
rect 49 -1044 51 -1034
rect 69 -1044 71 -1034
rect 151 -1068 153 -1058
rect 165 -1068 167 -1058
rect 185 -1068 187 -1058
rect 224 -1068 226 -1058
rect 238 -1068 240 -1058
rect 258 -1068 260 -1058
rect 296 -1070 298 -1060
rect 304 -1070 306 -1060
rect 321 -1070 323 -1060
rect 149 -1160 151 -1150
rect 163 -1160 165 -1150
rect 183 -1160 185 -1150
rect 215 -1162 217 -1152
rect 223 -1162 225 -1152
rect 240 -1162 242 -1152
rect 265 -1169 267 -1159
rect 273 -1169 275 -1159
rect 290 -1169 292 -1159
<< ptransistor >>
rect -3 -228 -1 -208
rect 11 -228 13 -208
rect 36 -219 38 -199
rect 50 -219 52 -199
rect 154 -221 156 -201
rect 168 -221 170 -201
rect 193 -212 195 -192
rect 207 -212 209 -192
rect 76 -242 78 -222
rect 90 -242 92 -222
rect 233 -235 235 -215
rect 247 -235 249 -215
rect 36 -288 38 -268
rect 50 -288 52 -268
rect 193 -281 195 -261
rect 207 -281 209 -261
rect 29 -354 31 -334
rect 43 -354 45 -334
rect 63 -354 65 -334
rect 145 -378 147 -358
rect 159 -378 161 -358
rect 179 -378 181 -358
rect 219 -383 221 -363
rect 226 -383 228 -363
rect 244 -383 246 -363
rect 3 -513 5 -493
rect 17 -513 19 -493
rect 42 -504 44 -484
rect 56 -504 58 -484
rect 160 -506 162 -486
rect 174 -506 176 -486
rect 199 -497 201 -477
rect 213 -497 215 -477
rect 82 -527 84 -507
rect 96 -527 98 -507
rect 239 -520 241 -500
rect 253 -520 255 -500
rect 42 -573 44 -553
rect 56 -573 58 -553
rect 199 -566 201 -546
rect 213 -566 215 -546
rect 35 -639 37 -619
rect 49 -639 51 -619
rect 69 -639 71 -619
rect 151 -663 153 -643
rect 165 -663 167 -643
rect 185 -663 187 -643
rect 224 -663 226 -643
rect 238 -663 240 -643
rect 258 -663 260 -643
rect 295 -668 297 -648
rect 302 -668 304 -648
rect 320 -668 322 -648
rect 248 -749 250 -729
rect 255 -749 257 -729
rect 273 -749 275 -729
rect 3 -893 5 -873
rect 17 -893 19 -873
rect 42 -884 44 -864
rect 56 -884 58 -864
rect 160 -886 162 -866
rect 174 -886 176 -866
rect 199 -877 201 -857
rect 213 -877 215 -857
rect 82 -907 84 -887
rect 96 -907 98 -887
rect 239 -900 241 -880
rect 253 -900 255 -880
rect 42 -953 44 -933
rect 56 -953 58 -933
rect 199 -946 201 -926
rect 213 -946 215 -926
rect 35 -1019 37 -999
rect 49 -1019 51 -999
rect 69 -1019 71 -999
rect 151 -1043 153 -1023
rect 165 -1043 167 -1023
rect 185 -1043 187 -1023
rect 224 -1043 226 -1023
rect 238 -1043 240 -1023
rect 258 -1043 260 -1023
rect 296 -1048 298 -1028
rect 303 -1048 305 -1028
rect 321 -1048 323 -1028
rect 149 -1135 151 -1115
rect 163 -1135 165 -1115
rect 183 -1135 185 -1115
rect 215 -1140 217 -1120
rect 222 -1140 224 -1120
rect 240 -1140 242 -1120
rect 265 -1147 267 -1127
rect 272 -1147 274 -1127
rect 290 -1147 292 -1127
<< ndiffusion >>
rect -4 -253 -3 -243
rect -1 -253 11 -243
rect 13 -253 14 -243
rect 35 -244 36 -234
rect 38 -244 50 -234
rect 52 -244 53 -234
rect 153 -246 154 -236
rect 156 -246 168 -236
rect 170 -246 171 -236
rect 192 -237 193 -227
rect 195 -237 207 -227
rect 209 -237 210 -227
rect 75 -267 76 -257
rect 78 -267 90 -257
rect 92 -267 93 -257
rect 232 -260 233 -250
rect 235 -260 247 -250
rect 249 -260 250 -250
rect 35 -313 36 -303
rect 38 -313 50 -303
rect 52 -313 53 -303
rect 192 -306 193 -296
rect 195 -306 207 -296
rect 209 -306 210 -296
rect 28 -379 29 -369
rect 31 -379 43 -369
rect 45 -379 46 -369
rect 60 -379 63 -369
rect 65 -379 68 -369
rect 144 -403 145 -393
rect 147 -403 159 -393
rect 161 -403 162 -393
rect 176 -403 179 -393
rect 181 -403 184 -393
rect 217 -405 219 -395
rect 221 -405 222 -395
rect 226 -405 227 -395
rect 229 -405 231 -395
rect 243 -405 244 -395
rect 246 -405 247 -395
rect 2 -538 3 -528
rect 5 -538 17 -528
rect 19 -538 20 -528
rect 41 -529 42 -519
rect 44 -529 56 -519
rect 58 -529 59 -519
rect 159 -531 160 -521
rect 162 -531 174 -521
rect 176 -531 177 -521
rect 198 -522 199 -512
rect 201 -522 213 -512
rect 215 -522 216 -512
rect 81 -552 82 -542
rect 84 -552 96 -542
rect 98 -552 99 -542
rect 238 -545 239 -535
rect 241 -545 253 -535
rect 255 -545 256 -535
rect 41 -598 42 -588
rect 44 -598 56 -588
rect 58 -598 59 -588
rect 198 -591 199 -581
rect 201 -591 213 -581
rect 215 -591 216 -581
rect 34 -664 35 -654
rect 37 -664 49 -654
rect 51 -664 52 -654
rect 66 -664 69 -654
rect 71 -664 74 -654
rect 150 -688 151 -678
rect 153 -688 165 -678
rect 167 -688 168 -678
rect 182 -688 185 -678
rect 187 -688 190 -678
rect 223 -688 224 -678
rect 226 -688 238 -678
rect 240 -688 241 -678
rect 255 -688 258 -678
rect 260 -688 263 -678
rect 293 -690 295 -680
rect 297 -690 298 -680
rect 302 -690 303 -680
rect 305 -690 307 -680
rect 319 -690 320 -680
rect 322 -690 323 -680
rect 246 -771 248 -761
rect 250 -771 251 -761
rect 255 -771 256 -761
rect 258 -771 260 -761
rect 272 -771 273 -761
rect 275 -771 276 -761
rect 2 -918 3 -908
rect 5 -918 17 -908
rect 19 -918 20 -908
rect 41 -909 42 -899
rect 44 -909 56 -899
rect 58 -909 59 -899
rect 159 -911 160 -901
rect 162 -911 174 -901
rect 176 -911 177 -901
rect 198 -902 199 -892
rect 201 -902 213 -892
rect 215 -902 216 -892
rect 81 -932 82 -922
rect 84 -932 96 -922
rect 98 -932 99 -922
rect 238 -925 239 -915
rect 241 -925 253 -915
rect 255 -925 256 -915
rect 41 -978 42 -968
rect 44 -978 56 -968
rect 58 -978 59 -968
rect 198 -971 199 -961
rect 201 -971 213 -961
rect 215 -971 216 -961
rect 34 -1044 35 -1034
rect 37 -1044 49 -1034
rect 51 -1044 52 -1034
rect 66 -1044 69 -1034
rect 71 -1044 74 -1034
rect 150 -1068 151 -1058
rect 153 -1068 165 -1058
rect 167 -1068 168 -1058
rect 182 -1068 185 -1058
rect 187 -1068 190 -1058
rect 223 -1068 224 -1058
rect 226 -1068 238 -1058
rect 240 -1068 241 -1058
rect 255 -1068 258 -1058
rect 260 -1068 263 -1058
rect 294 -1070 296 -1060
rect 298 -1070 299 -1060
rect 303 -1070 304 -1060
rect 306 -1070 308 -1060
rect 320 -1070 321 -1060
rect 323 -1070 324 -1060
rect 148 -1160 149 -1150
rect 151 -1160 163 -1150
rect 165 -1160 166 -1150
rect 180 -1160 183 -1150
rect 185 -1160 188 -1150
rect 213 -1162 215 -1152
rect 217 -1162 218 -1152
rect 222 -1162 223 -1152
rect 225 -1162 227 -1152
rect 239 -1162 240 -1152
rect 242 -1162 243 -1152
rect 263 -1169 265 -1159
rect 267 -1169 268 -1159
rect 272 -1169 273 -1159
rect 275 -1169 277 -1159
rect 289 -1169 290 -1159
rect 292 -1169 293 -1159
<< pdiffusion >>
rect -4 -228 -3 -208
rect -1 -228 3 -208
rect 7 -228 11 -208
rect 13 -228 14 -208
rect 35 -219 36 -199
rect 38 -219 42 -199
rect 46 -219 50 -199
rect 52 -219 53 -199
rect 153 -221 154 -201
rect 156 -221 160 -201
rect 164 -221 168 -201
rect 170 -221 171 -201
rect 192 -212 193 -192
rect 195 -212 199 -192
rect 203 -212 207 -192
rect 209 -212 210 -192
rect 75 -242 76 -222
rect 78 -242 82 -222
rect 86 -242 90 -222
rect 92 -242 93 -222
rect 232 -235 233 -215
rect 235 -235 239 -215
rect 243 -235 247 -215
rect 249 -235 250 -215
rect 35 -288 36 -268
rect 38 -288 42 -268
rect 46 -288 50 -268
rect 52 -288 53 -268
rect 192 -281 193 -261
rect 195 -281 199 -261
rect 203 -281 207 -261
rect 209 -281 210 -261
rect 28 -354 29 -334
rect 31 -354 35 -334
rect 39 -354 43 -334
rect 45 -354 46 -334
rect 60 -354 63 -334
rect 65 -354 68 -334
rect 144 -378 145 -358
rect 147 -378 151 -358
rect 155 -378 159 -358
rect 161 -378 162 -358
rect 176 -378 179 -358
rect 181 -378 184 -358
rect 217 -383 219 -363
rect 221 -383 226 -363
rect 228 -383 230 -363
rect 243 -383 244 -363
rect 246 -383 247 -363
rect 2 -513 3 -493
rect 5 -513 9 -493
rect 13 -513 17 -493
rect 19 -513 20 -493
rect 41 -504 42 -484
rect 44 -504 48 -484
rect 52 -504 56 -484
rect 58 -504 59 -484
rect 159 -506 160 -486
rect 162 -506 166 -486
rect 170 -506 174 -486
rect 176 -506 177 -486
rect 198 -497 199 -477
rect 201 -497 205 -477
rect 209 -497 213 -477
rect 215 -497 216 -477
rect 81 -527 82 -507
rect 84 -527 88 -507
rect 92 -527 96 -507
rect 98 -527 99 -507
rect 238 -520 239 -500
rect 241 -520 245 -500
rect 249 -520 253 -500
rect 255 -520 256 -500
rect 41 -573 42 -553
rect 44 -573 48 -553
rect 52 -573 56 -553
rect 58 -573 59 -553
rect 198 -566 199 -546
rect 201 -566 205 -546
rect 209 -566 213 -546
rect 215 -566 216 -546
rect 34 -639 35 -619
rect 37 -639 41 -619
rect 45 -639 49 -619
rect 51 -639 52 -619
rect 66 -639 69 -619
rect 71 -639 74 -619
rect 150 -663 151 -643
rect 153 -663 157 -643
rect 161 -663 165 -643
rect 167 -663 168 -643
rect 182 -663 185 -643
rect 187 -663 190 -643
rect 223 -663 224 -643
rect 226 -663 230 -643
rect 234 -663 238 -643
rect 240 -663 241 -643
rect 255 -663 258 -643
rect 260 -663 263 -643
rect 293 -668 295 -648
rect 297 -668 302 -648
rect 304 -668 306 -648
rect 319 -668 320 -648
rect 322 -668 323 -648
rect 246 -749 248 -729
rect 250 -749 255 -729
rect 257 -749 259 -729
rect 272 -749 273 -729
rect 275 -749 276 -729
rect 2 -893 3 -873
rect 5 -893 9 -873
rect 13 -893 17 -873
rect 19 -893 20 -873
rect 41 -884 42 -864
rect 44 -884 48 -864
rect 52 -884 56 -864
rect 58 -884 59 -864
rect 159 -886 160 -866
rect 162 -886 166 -866
rect 170 -886 174 -866
rect 176 -886 177 -866
rect 198 -877 199 -857
rect 201 -877 205 -857
rect 209 -877 213 -857
rect 215 -877 216 -857
rect 81 -907 82 -887
rect 84 -907 88 -887
rect 92 -907 96 -887
rect 98 -907 99 -887
rect 238 -900 239 -880
rect 241 -900 245 -880
rect 249 -900 253 -880
rect 255 -900 256 -880
rect 41 -953 42 -933
rect 44 -953 48 -933
rect 52 -953 56 -933
rect 58 -953 59 -933
rect 198 -946 199 -926
rect 201 -946 205 -926
rect 209 -946 213 -926
rect 215 -946 216 -926
rect 34 -1019 35 -999
rect 37 -1019 41 -999
rect 45 -1019 49 -999
rect 51 -1019 52 -999
rect 66 -1019 69 -999
rect 71 -1019 74 -999
rect 150 -1043 151 -1023
rect 153 -1043 157 -1023
rect 161 -1043 165 -1023
rect 167 -1043 168 -1023
rect 182 -1043 185 -1023
rect 187 -1043 190 -1023
rect 223 -1043 224 -1023
rect 226 -1043 230 -1023
rect 234 -1043 238 -1023
rect 240 -1043 241 -1023
rect 255 -1043 258 -1023
rect 260 -1043 263 -1023
rect 294 -1048 296 -1028
rect 298 -1048 303 -1028
rect 305 -1048 307 -1028
rect 320 -1048 321 -1028
rect 323 -1048 324 -1028
rect 148 -1135 149 -1115
rect 151 -1135 155 -1115
rect 159 -1135 163 -1115
rect 165 -1135 166 -1115
rect 180 -1135 183 -1115
rect 185 -1135 188 -1115
rect 213 -1140 215 -1120
rect 217 -1140 222 -1120
rect 224 -1140 226 -1120
rect 239 -1140 240 -1120
rect 242 -1140 243 -1120
rect 263 -1147 265 -1127
rect 267 -1147 272 -1127
rect 274 -1147 276 -1127
rect 289 -1147 290 -1127
rect 292 -1147 293 -1127
<< ndcontact >>
rect -8 -253 -4 -243
rect 14 -253 18 -243
rect 31 -244 35 -234
rect 53 -244 57 -234
rect 149 -246 153 -236
rect 171 -246 175 -236
rect 188 -237 192 -227
rect 210 -237 214 -227
rect 71 -267 75 -257
rect 93 -267 97 -257
rect 228 -260 232 -250
rect 250 -260 254 -250
rect 31 -313 35 -303
rect 53 -313 57 -303
rect 188 -306 192 -296
rect 210 -306 214 -296
rect 24 -379 28 -369
rect 46 -379 50 -369
rect 56 -379 60 -369
rect 68 -379 72 -369
rect 140 -403 144 -393
rect 162 -403 166 -393
rect 172 -403 176 -393
rect 184 -403 188 -393
rect 213 -405 217 -395
rect 222 -405 226 -395
rect 231 -405 235 -395
rect 239 -405 243 -395
rect 247 -405 251 -395
rect -2 -538 2 -528
rect 20 -538 24 -528
rect 37 -529 41 -519
rect 59 -529 63 -519
rect 155 -531 159 -521
rect 177 -531 181 -521
rect 194 -522 198 -512
rect 216 -522 220 -512
rect 77 -552 81 -542
rect 99 -552 103 -542
rect 234 -545 238 -535
rect 256 -545 260 -535
rect 37 -598 41 -588
rect 59 -598 63 -588
rect 194 -591 198 -581
rect 216 -591 220 -581
rect 30 -664 34 -654
rect 52 -664 56 -654
rect 62 -664 66 -654
rect 74 -664 78 -654
rect 146 -688 150 -678
rect 168 -688 172 -678
rect 178 -688 182 -678
rect 190 -688 194 -678
rect 219 -688 223 -678
rect 241 -688 245 -678
rect 251 -688 255 -678
rect 263 -688 267 -678
rect 289 -690 293 -680
rect 298 -690 302 -680
rect 307 -690 311 -680
rect 315 -690 319 -680
rect 323 -690 327 -680
rect 242 -771 246 -761
rect 251 -771 255 -761
rect 260 -771 264 -761
rect 268 -771 272 -761
rect 276 -771 280 -761
rect -2 -918 2 -908
rect 20 -918 24 -908
rect 37 -909 41 -899
rect 59 -909 63 -899
rect 155 -911 159 -901
rect 177 -911 181 -901
rect 194 -902 198 -892
rect 216 -902 220 -892
rect 77 -932 81 -922
rect 99 -932 103 -922
rect 234 -925 238 -915
rect 256 -925 260 -915
rect 37 -978 41 -968
rect 59 -978 63 -968
rect 194 -971 198 -961
rect 216 -971 220 -961
rect 30 -1044 34 -1034
rect 52 -1044 56 -1034
rect 62 -1044 66 -1034
rect 74 -1044 78 -1034
rect 146 -1068 150 -1058
rect 168 -1068 172 -1058
rect 178 -1068 182 -1058
rect 190 -1068 194 -1058
rect 219 -1068 223 -1058
rect 241 -1068 245 -1058
rect 251 -1068 255 -1058
rect 263 -1068 267 -1058
rect 290 -1070 294 -1060
rect 299 -1070 303 -1060
rect 308 -1070 312 -1060
rect 316 -1070 320 -1060
rect 324 -1070 328 -1060
rect 144 -1160 148 -1150
rect 166 -1160 170 -1150
rect 176 -1160 180 -1150
rect 188 -1160 192 -1150
rect 209 -1162 213 -1152
rect 218 -1162 222 -1152
rect 227 -1162 231 -1152
rect 235 -1162 239 -1152
rect 243 -1162 247 -1152
rect 259 -1169 263 -1159
rect 268 -1169 272 -1159
rect 277 -1169 281 -1159
rect 285 -1169 289 -1159
rect 293 -1169 297 -1159
<< pdcontact >>
rect -8 -228 -4 -208
rect 3 -228 7 -208
rect 14 -228 18 -208
rect 31 -219 35 -199
rect 42 -219 46 -199
rect 53 -219 57 -199
rect 149 -221 153 -201
rect 160 -221 164 -201
rect 171 -221 175 -201
rect 188 -212 192 -192
rect 199 -212 203 -192
rect 210 -212 214 -192
rect 71 -242 75 -222
rect 82 -242 86 -222
rect 93 -242 97 -222
rect 228 -235 232 -215
rect 239 -235 243 -215
rect 250 -235 254 -215
rect 31 -288 35 -268
rect 42 -288 46 -268
rect 53 -288 57 -268
rect 188 -281 192 -261
rect 199 -281 203 -261
rect 210 -281 214 -261
rect 24 -354 28 -334
rect 35 -354 39 -334
rect 46 -354 50 -334
rect 56 -354 60 -334
rect 68 -354 72 -334
rect 140 -378 144 -358
rect 151 -378 155 -358
rect 162 -378 166 -358
rect 172 -378 176 -358
rect 184 -378 188 -358
rect 213 -383 217 -363
rect 230 -383 234 -363
rect 239 -383 243 -363
rect 247 -383 251 -363
rect -2 -513 2 -493
rect 9 -513 13 -493
rect 20 -513 24 -493
rect 37 -504 41 -484
rect 48 -504 52 -484
rect 59 -504 63 -484
rect 155 -506 159 -486
rect 166 -506 170 -486
rect 177 -506 181 -486
rect 194 -497 198 -477
rect 205 -497 209 -477
rect 216 -497 220 -477
rect 77 -527 81 -507
rect 88 -527 92 -507
rect 99 -527 103 -507
rect 234 -520 238 -500
rect 245 -520 249 -500
rect 256 -520 260 -500
rect 37 -573 41 -553
rect 48 -573 52 -553
rect 59 -573 63 -553
rect 194 -566 198 -546
rect 205 -566 209 -546
rect 216 -566 220 -546
rect 30 -639 34 -619
rect 41 -639 45 -619
rect 52 -639 56 -619
rect 62 -639 66 -619
rect 74 -639 78 -619
rect 146 -663 150 -643
rect 157 -663 161 -643
rect 168 -663 172 -643
rect 178 -663 182 -643
rect 190 -663 194 -643
rect 219 -663 223 -643
rect 230 -663 234 -643
rect 241 -663 245 -643
rect 251 -663 255 -643
rect 263 -663 267 -643
rect 289 -668 293 -648
rect 306 -668 310 -648
rect 315 -668 319 -648
rect 323 -668 327 -648
rect 242 -749 246 -729
rect 259 -749 263 -729
rect 268 -749 272 -729
rect 276 -749 280 -729
rect -2 -893 2 -873
rect 9 -893 13 -873
rect 20 -893 24 -873
rect 37 -884 41 -864
rect 48 -884 52 -864
rect 59 -884 63 -864
rect 155 -886 159 -866
rect 166 -886 170 -866
rect 177 -886 181 -866
rect 194 -877 198 -857
rect 205 -877 209 -857
rect 216 -877 220 -857
rect 77 -907 81 -887
rect 88 -907 92 -887
rect 99 -907 103 -887
rect 234 -900 238 -880
rect 245 -900 249 -880
rect 256 -900 260 -880
rect 37 -953 41 -933
rect 48 -953 52 -933
rect 59 -953 63 -933
rect 194 -946 198 -926
rect 205 -946 209 -926
rect 216 -946 220 -926
rect 30 -1019 34 -999
rect 41 -1019 45 -999
rect 52 -1019 56 -999
rect 62 -1019 66 -999
rect 74 -1019 78 -999
rect 146 -1043 150 -1023
rect 157 -1043 161 -1023
rect 168 -1043 172 -1023
rect 178 -1043 182 -1023
rect 190 -1043 194 -1023
rect 219 -1043 223 -1023
rect 230 -1043 234 -1023
rect 241 -1043 245 -1023
rect 251 -1043 255 -1023
rect 263 -1043 267 -1023
rect 290 -1048 294 -1028
rect 307 -1048 311 -1028
rect 316 -1048 320 -1028
rect 324 -1048 328 -1028
rect 144 -1135 148 -1115
rect 155 -1135 159 -1115
rect 166 -1135 170 -1115
rect 176 -1135 180 -1115
rect 188 -1135 192 -1115
rect 209 -1140 213 -1120
rect 226 -1140 230 -1120
rect 235 -1140 239 -1120
rect 243 -1140 247 -1120
rect 259 -1147 263 -1127
rect 276 -1147 280 -1127
rect 285 -1147 289 -1127
rect 293 -1147 297 -1127
<< polysilicon >>
rect 98 -77 100 -76
rect 105 -77 107 -76
rect 193 -192 195 -189
rect 207 -192 209 -189
rect 36 -199 38 -196
rect 50 -199 52 -196
rect -3 -208 -1 -205
rect 11 -208 13 -205
rect 154 -201 156 -198
rect 168 -201 170 -198
rect -3 -243 -1 -228
rect 11 -243 13 -228
rect 36 -234 38 -219
rect 50 -234 52 -219
rect 76 -222 78 -219
rect 90 -222 92 -219
rect 154 -236 156 -221
rect 168 -236 170 -221
rect 193 -227 195 -212
rect 207 -227 209 -212
rect 233 -215 235 -212
rect 247 -215 249 -212
rect 36 -249 38 -244
rect 50 -249 52 -244
rect -3 -258 -1 -253
rect 11 -258 13 -253
rect 76 -257 78 -242
rect 90 -257 92 -242
rect 193 -242 195 -237
rect 207 -242 209 -237
rect 154 -251 156 -246
rect 168 -251 170 -246
rect 233 -250 235 -235
rect 247 -250 249 -235
rect 36 -268 38 -265
rect 50 -268 52 -265
rect 193 -261 195 -258
rect 207 -261 209 -258
rect 76 -272 78 -267
rect 90 -272 92 -267
rect 233 -265 235 -260
rect 247 -265 249 -260
rect 36 -303 38 -288
rect 50 -303 52 -288
rect 193 -296 195 -281
rect 207 -296 209 -281
rect 193 -311 195 -306
rect 207 -311 209 -306
rect 36 -318 38 -313
rect 50 -318 52 -313
rect 29 -334 31 -331
rect 43 -334 45 -331
rect 63 -334 65 -331
rect 29 -369 31 -354
rect 43 -369 45 -354
rect 63 -369 65 -354
rect 145 -358 147 -355
rect 159 -358 161 -355
rect 179 -358 181 -355
rect 219 -363 221 -349
rect 226 -363 228 -349
rect 244 -363 246 -360
rect 29 -384 31 -379
rect 43 -384 45 -379
rect 63 -382 65 -379
rect 145 -393 147 -378
rect 159 -393 161 -378
rect 179 -393 181 -378
rect 219 -395 221 -383
rect 226 -391 228 -383
rect 226 -393 229 -391
rect 227 -395 229 -393
rect 244 -395 246 -383
rect 145 -408 147 -403
rect 159 -408 161 -403
rect 179 -406 181 -403
rect 219 -408 221 -405
rect 227 -408 229 -405
rect 244 -408 246 -405
rect 199 -477 201 -474
rect 213 -477 215 -474
rect 42 -484 44 -481
rect 56 -484 58 -481
rect 3 -493 5 -490
rect 17 -493 19 -490
rect 160 -486 162 -483
rect 174 -486 176 -483
rect 3 -528 5 -513
rect 17 -528 19 -513
rect 42 -519 44 -504
rect 56 -519 58 -504
rect 82 -507 84 -504
rect 96 -507 98 -504
rect 160 -521 162 -506
rect 174 -521 176 -506
rect 199 -512 201 -497
rect 213 -512 215 -497
rect 239 -500 241 -497
rect 253 -500 255 -497
rect 42 -534 44 -529
rect 56 -534 58 -529
rect 3 -543 5 -538
rect 17 -543 19 -538
rect 82 -542 84 -527
rect 96 -542 98 -527
rect 199 -527 201 -522
rect 213 -527 215 -522
rect 160 -536 162 -531
rect 174 -536 176 -531
rect 239 -535 241 -520
rect 253 -535 255 -520
rect 42 -553 44 -550
rect 56 -553 58 -550
rect 199 -546 201 -543
rect 213 -546 215 -543
rect 82 -557 84 -552
rect 96 -557 98 -552
rect 239 -550 241 -545
rect 253 -550 255 -545
rect 42 -588 44 -573
rect 56 -588 58 -573
rect 199 -581 201 -566
rect 213 -581 215 -566
rect 199 -596 201 -591
rect 213 -596 215 -591
rect 42 -603 44 -598
rect 56 -603 58 -598
rect 35 -619 37 -616
rect 49 -619 51 -616
rect 69 -619 71 -616
rect 35 -654 37 -639
rect 49 -654 51 -639
rect 69 -654 71 -639
rect 151 -643 153 -640
rect 165 -643 167 -640
rect 185 -643 187 -640
rect 224 -643 226 -640
rect 238 -643 240 -640
rect 258 -643 260 -640
rect 295 -648 297 -634
rect 302 -648 304 -634
rect 320 -648 322 -645
rect 35 -669 37 -664
rect 49 -669 51 -664
rect 69 -667 71 -664
rect 151 -678 153 -663
rect 165 -678 167 -663
rect 185 -678 187 -663
rect 224 -678 226 -663
rect 238 -678 240 -663
rect 258 -678 260 -663
rect 295 -680 297 -668
rect 302 -676 304 -668
rect 302 -678 305 -676
rect 303 -680 305 -678
rect 320 -680 322 -668
rect 151 -693 153 -688
rect 165 -693 167 -688
rect 185 -691 187 -688
rect 224 -693 226 -688
rect 238 -693 240 -688
rect 258 -691 260 -688
rect 295 -693 297 -690
rect 303 -693 305 -690
rect 320 -693 322 -690
rect 248 -729 250 -715
rect 255 -729 257 -715
rect 273 -729 275 -726
rect 248 -761 250 -749
rect 255 -757 257 -749
rect 255 -759 258 -757
rect 256 -761 258 -759
rect 273 -761 275 -749
rect 248 -774 250 -771
rect 256 -774 258 -771
rect 273 -774 275 -771
rect 199 -857 201 -854
rect 213 -857 215 -854
rect 42 -864 44 -861
rect 56 -864 58 -861
rect 3 -873 5 -870
rect 17 -873 19 -870
rect 160 -866 162 -863
rect 174 -866 176 -863
rect 3 -908 5 -893
rect 17 -908 19 -893
rect 42 -899 44 -884
rect 56 -899 58 -884
rect 82 -887 84 -884
rect 96 -887 98 -884
rect 160 -901 162 -886
rect 174 -901 176 -886
rect 199 -892 201 -877
rect 213 -892 215 -877
rect 239 -880 241 -877
rect 253 -880 255 -877
rect 42 -914 44 -909
rect 56 -914 58 -909
rect 3 -923 5 -918
rect 17 -923 19 -918
rect 82 -922 84 -907
rect 96 -922 98 -907
rect 199 -906 201 -902
rect 213 -907 215 -902
rect 160 -916 162 -911
rect 174 -916 176 -911
rect 239 -915 241 -900
rect 253 -915 255 -900
rect 42 -933 44 -930
rect 56 -933 58 -930
rect 199 -926 201 -923
rect 213 -926 215 -923
rect 82 -937 84 -932
rect 96 -937 98 -932
rect 239 -930 241 -925
rect 253 -930 255 -925
rect 42 -968 44 -953
rect 56 -968 58 -953
rect 199 -961 201 -946
rect 213 -961 215 -946
rect 199 -976 201 -971
rect 213 -976 215 -971
rect 42 -983 44 -978
rect 56 -983 58 -978
rect 35 -999 37 -996
rect 49 -999 51 -996
rect 69 -999 71 -996
rect 35 -1034 37 -1019
rect 49 -1034 51 -1019
rect 69 -1034 71 -1019
rect 151 -1023 153 -1020
rect 165 -1023 167 -1020
rect 185 -1023 187 -1020
rect 224 -1023 226 -1020
rect 238 -1023 240 -1020
rect 258 -1023 260 -1020
rect 296 -1028 298 -1014
rect 303 -1028 305 -1014
rect 321 -1028 323 -1025
rect 35 -1049 37 -1044
rect 49 -1049 51 -1044
rect 69 -1047 71 -1044
rect 151 -1058 153 -1043
rect 165 -1058 167 -1043
rect 185 -1058 187 -1043
rect 224 -1058 226 -1043
rect 238 -1058 240 -1043
rect 258 -1058 260 -1043
rect 296 -1060 298 -1048
rect 303 -1056 305 -1048
rect 303 -1058 306 -1056
rect 304 -1060 306 -1058
rect 321 -1060 323 -1048
rect 151 -1073 153 -1068
rect 165 -1073 167 -1068
rect 185 -1071 187 -1068
rect 224 -1073 226 -1068
rect 238 -1073 240 -1068
rect 258 -1071 260 -1068
rect 296 -1073 298 -1070
rect 304 -1073 306 -1070
rect 321 -1073 323 -1070
rect 149 -1115 151 -1112
rect 163 -1115 165 -1112
rect 183 -1115 185 -1112
rect 215 -1120 217 -1106
rect 222 -1120 224 -1106
rect 240 -1120 242 -1117
rect 149 -1150 151 -1135
rect 163 -1150 165 -1135
rect 183 -1150 185 -1135
rect 265 -1127 267 -1113
rect 272 -1127 274 -1113
rect 290 -1127 292 -1124
rect 215 -1152 217 -1140
rect 222 -1148 224 -1140
rect 222 -1150 225 -1148
rect 223 -1152 225 -1150
rect 240 -1152 242 -1140
rect 149 -1165 151 -1160
rect 163 -1165 165 -1160
rect 183 -1163 185 -1160
rect 265 -1159 267 -1147
rect 272 -1155 274 -1147
rect 272 -1157 275 -1155
rect 273 -1159 275 -1157
rect 290 -1159 292 -1147
rect 215 -1165 217 -1162
rect 223 -1165 225 -1162
rect 240 -1165 242 -1162
rect 265 -1172 267 -1169
rect 273 -1172 275 -1169
rect 290 -1172 292 -1169
<< polycontact >>
rect 94 -80 98 -76
rect 107 -80 111 -76
rect 32 -230 36 -226
rect 189 -223 193 -219
rect 46 -249 50 -245
rect 72 -251 76 -247
rect -1 -258 3 -254
rect 7 -258 11 -254
rect 86 -256 90 -252
rect 203 -242 207 -238
rect 229 -244 233 -240
rect 156 -251 160 -247
rect 164 -251 168 -247
rect 243 -249 247 -245
rect 32 -297 36 -293
rect 189 -290 193 -286
rect 203 -311 207 -307
rect 46 -318 50 -314
rect 215 -353 219 -349
rect 25 -366 29 -362
rect 39 -368 43 -364
rect 59 -361 63 -357
rect 228 -353 232 -349
rect 141 -390 145 -386
rect 155 -392 159 -388
rect 175 -385 179 -381
rect 240 -390 244 -386
rect 38 -515 42 -511
rect 195 -508 199 -504
rect 52 -534 56 -530
rect 78 -536 82 -532
rect 5 -543 9 -539
rect 13 -543 17 -539
rect 92 -541 96 -537
rect 209 -527 213 -523
rect 235 -529 239 -525
rect 162 -536 166 -532
rect 170 -536 174 -532
rect 249 -534 253 -530
rect 38 -582 42 -578
rect 195 -575 199 -571
rect 209 -596 213 -592
rect 52 -603 56 -599
rect 291 -638 295 -634
rect 31 -651 35 -647
rect 45 -653 49 -649
rect 65 -646 69 -642
rect 304 -638 308 -634
rect 147 -675 151 -671
rect 161 -677 165 -673
rect 181 -670 185 -666
rect 220 -675 224 -671
rect 234 -677 238 -673
rect 254 -670 258 -666
rect 316 -675 320 -671
rect 244 -719 248 -715
rect 257 -719 261 -715
rect 269 -756 273 -752
rect 38 -895 42 -891
rect 195 -888 199 -884
rect 52 -914 56 -910
rect 78 -916 82 -912
rect 5 -923 9 -919
rect 13 -923 17 -919
rect 92 -921 96 -917
rect 209 -907 213 -903
rect 235 -909 239 -905
rect 162 -916 166 -912
rect 170 -916 174 -912
rect 249 -914 253 -910
rect 38 -962 42 -958
rect 195 -955 199 -951
rect 209 -976 213 -972
rect 52 -983 56 -979
rect 292 -1018 296 -1014
rect 31 -1031 35 -1027
rect 45 -1033 49 -1029
rect 65 -1026 69 -1022
rect 305 -1018 309 -1014
rect 147 -1055 151 -1051
rect 161 -1057 165 -1053
rect 181 -1050 185 -1046
rect 220 -1055 224 -1051
rect 234 -1057 238 -1053
rect 254 -1050 258 -1046
rect 317 -1055 321 -1051
rect 211 -1110 215 -1106
rect 224 -1110 228 -1106
rect 261 -1117 265 -1113
rect 145 -1147 149 -1143
rect 159 -1149 163 -1145
rect 179 -1142 183 -1138
rect 274 -1117 278 -1113
rect 236 -1147 240 -1143
rect 286 -1154 290 -1150
<< metal1 >>
rect 229 65 234 67
rect 39 58 43 62
rect 103 50 174 53
rect -43 34 -20 37
rect -43 25 -29 28
rect -32 -22 -29 25
rect -23 -14 -20 34
rect 103 4 106 50
rect 123 45 128 47
rect 111 34 115 37
rect 45 0 47 4
rect 103 2 113 4
rect 105 0 113 2
rect 110 -3 113 0
rect -13 -10 -7 -7
rect 30 -8 36 -6
rect -13 -13 -11 -10
rect 0 -16 4 -9
rect -18 -19 4 -16
rect 8 -22 12 -9
rect 47 -12 53 -9
rect -32 -25 12 -22
rect -32 -144 -29 -25
rect 67 -29 76 -27
rect 131 -29 138 -25
rect -23 -114 -20 -36
rect 45 -69 47 -65
rect 45 -77 48 -75
rect 165 -76 168 6
rect 171 -9 174 50
rect 234 7 236 11
rect 287 6 289 7
rect 225 1 227 5
rect 178 -2 183 0
rect 235 -2 241 -1
rect 189 -9 193 -2
rect 171 -13 193 -9
rect 179 -14 182 -13
rect 197 -73 201 -2
rect 234 -5 241 -2
rect 256 -22 265 -20
rect 214 -66 217 -62
rect 236 -64 240 -62
rect 311 -64 314 77
rect 323 7 326 10
rect 236 -67 314 -64
rect 236 -73 240 -67
rect 197 -76 240 -73
rect 78 -80 94 -76
rect 111 -80 168 -76
rect 78 -108 81 -80
rect 89 -87 91 -83
rect 76 -112 81 -108
rect -23 -117 24 -114
rect 51 -142 57 -139
rect 29 -144 35 -142
rect -32 -147 35 -144
rect 78 -162 81 -112
rect 131 -116 281 -113
rect 105 -142 108 -139
rect 78 -166 202 -162
rect 171 -188 232 -184
rect 14 -195 75 -191
rect 171 -193 175 -188
rect 14 -200 18 -195
rect -12 -204 18 -200
rect -8 -208 -4 -204
rect 14 -208 18 -204
rect -44 -215 -21 -212
rect -44 -224 -30 -221
rect -33 -271 -30 -224
rect -24 -263 -21 -215
rect 31 -199 35 -195
rect 53 -199 57 -195
rect 71 -214 75 -195
rect 149 -197 175 -193
rect 149 -201 153 -197
rect 171 -201 175 -197
rect 71 -218 97 -214
rect 42 -222 46 -219
rect 71 -222 75 -218
rect 93 -222 97 -218
rect 188 -192 192 -188
rect 210 -192 214 -188
rect 228 -207 232 -188
rect 228 -211 254 -207
rect 199 -215 203 -212
rect 228 -215 232 -211
rect 250 -215 254 -211
rect 199 -219 221 -215
rect 42 -226 64 -222
rect 3 -231 7 -228
rect 22 -230 32 -226
rect 22 -231 26 -230
rect 3 -235 26 -231
rect 53 -234 57 -226
rect 14 -243 18 -235
rect -8 -258 -4 -253
rect -12 -262 -4 -258
rect -1 -265 3 -258
rect -19 -268 3 -265
rect 7 -271 11 -258
rect -33 -274 11 -271
rect -33 -393 -30 -274
rect -24 -363 -21 -285
rect 22 -293 26 -235
rect 31 -249 35 -244
rect 44 -249 46 -245
rect 60 -247 64 -226
rect 160 -224 164 -221
rect 179 -223 189 -219
rect 179 -224 183 -223
rect 160 -228 183 -224
rect 210 -227 214 -219
rect 171 -236 175 -228
rect 82 -245 86 -242
rect 29 -255 35 -249
rect 60 -251 72 -247
rect 82 -249 141 -245
rect 81 -256 86 -252
rect 42 -260 46 -257
rect 31 -264 57 -260
rect 31 -268 35 -264
rect 53 -268 57 -264
rect 71 -272 75 -267
rect 66 -276 75 -272
rect 42 -291 46 -288
rect 81 -291 85 -256
rect 93 -257 97 -249
rect 22 -297 32 -293
rect 42 -295 85 -291
rect 53 -303 57 -295
rect 31 -318 35 -313
rect 44 -318 46 -314
rect 26 -322 35 -318
rect 24 -329 60 -326
rect 24 -330 50 -329
rect 24 -334 28 -330
rect 46 -334 50 -330
rect 56 -334 60 -329
rect 35 -357 39 -354
rect 68 -357 72 -354
rect 35 -361 59 -357
rect 68 -361 96 -357
rect 23 -363 25 -362
rect -24 -366 25 -363
rect 46 -369 50 -361
rect 68 -369 72 -361
rect 24 -384 28 -379
rect 22 -385 28 -384
rect 56 -385 60 -379
rect 22 -388 60 -385
rect 28 -393 34 -391
rect -33 -396 34 -393
rect 92 -430 96 -361
rect 131 -386 134 -249
rect 138 -258 141 -249
rect 149 -251 153 -246
rect 145 -255 153 -251
rect 156 -258 160 -251
rect 138 -262 160 -258
rect 164 -322 167 -251
rect 179 -286 183 -228
rect 188 -242 192 -237
rect 201 -242 203 -238
rect 217 -240 221 -219
rect 239 -238 243 -235
rect 186 -248 192 -242
rect 217 -244 229 -240
rect 239 -242 256 -238
rect 250 -243 256 -242
rect 238 -249 243 -245
rect 199 -253 203 -250
rect 188 -257 214 -253
rect 188 -261 192 -257
rect 210 -261 214 -257
rect 228 -265 232 -260
rect 223 -269 232 -265
rect 199 -284 203 -281
rect 238 -284 242 -249
rect 250 -250 254 -243
rect 179 -290 189 -286
rect 199 -288 242 -284
rect 210 -296 214 -288
rect 188 -311 192 -306
rect 183 -315 192 -311
rect 203 -313 207 -311
rect 278 -313 281 -116
rect 303 -165 372 -162
rect 290 -242 292 -239
rect 203 -316 281 -313
rect 203 -322 206 -316
rect 164 -325 206 -322
rect 369 -338 372 -165
rect 149 -341 372 -338
rect 149 -342 154 -341
rect 369 -343 372 -341
rect 140 -353 176 -350
rect 140 -354 166 -353
rect 140 -358 144 -354
rect 162 -358 166 -354
rect 172 -358 176 -353
rect 191 -353 215 -349
rect 232 -353 269 -349
rect 151 -381 155 -378
rect 184 -381 188 -378
rect 191 -380 194 -353
rect 210 -359 243 -356
rect 210 -360 217 -359
rect 213 -363 217 -360
rect 239 -363 243 -359
rect 151 -385 175 -381
rect 184 -385 191 -381
rect 131 -390 141 -386
rect 154 -392 155 -388
rect 162 -393 166 -385
rect 184 -393 188 -385
rect 230 -386 234 -383
rect 247 -386 251 -383
rect 222 -390 240 -386
rect 247 -389 255 -386
rect 222 -395 226 -390
rect 247 -395 251 -389
rect 140 -409 144 -403
rect 172 -409 176 -403
rect 140 -412 176 -409
rect 213 -409 217 -405
rect 231 -409 235 -405
rect 239 -409 243 -405
rect 213 -412 243 -409
rect 157 -416 164 -412
rect 226 -415 229 -412
rect 266 -430 269 -353
rect 92 -433 362 -430
rect 256 -456 259 -443
rect 256 -459 287 -456
rect 177 -473 238 -469
rect 20 -480 81 -476
rect 177 -478 181 -473
rect 20 -485 24 -480
rect -6 -489 24 -485
rect -2 -493 2 -489
rect 20 -493 24 -489
rect -38 -500 -15 -497
rect -38 -509 -24 -506
rect -27 -556 -24 -509
rect -18 -548 -15 -500
rect 37 -484 41 -480
rect 59 -484 63 -480
rect 77 -499 81 -480
rect 155 -482 181 -478
rect 155 -486 159 -482
rect 177 -486 181 -482
rect 77 -503 103 -499
rect 48 -507 52 -504
rect 77 -507 81 -503
rect 99 -507 103 -503
rect 194 -477 198 -473
rect 216 -477 220 -473
rect 234 -492 238 -473
rect 234 -496 260 -492
rect 205 -500 209 -497
rect 234 -500 238 -496
rect 256 -500 260 -496
rect 205 -504 227 -500
rect 48 -511 70 -507
rect 9 -516 13 -513
rect 28 -515 38 -511
rect 28 -516 32 -515
rect 9 -520 32 -516
rect 59 -519 63 -511
rect 20 -528 24 -520
rect -2 -543 2 -538
rect -6 -547 2 -543
rect 5 -550 9 -543
rect -13 -553 9 -550
rect 13 -556 17 -543
rect -27 -559 17 -556
rect -27 -678 -24 -559
rect -18 -648 -15 -570
rect 28 -578 32 -520
rect 37 -534 41 -529
rect 50 -534 52 -530
rect 66 -532 70 -511
rect 166 -509 170 -506
rect 185 -508 195 -504
rect 185 -509 189 -508
rect 166 -513 189 -509
rect 216 -512 220 -504
rect 177 -521 181 -513
rect 88 -530 92 -527
rect 35 -540 41 -534
rect 66 -536 78 -532
rect 88 -534 147 -530
rect 87 -541 92 -537
rect 48 -545 52 -542
rect 37 -549 63 -545
rect 37 -553 41 -549
rect 59 -553 63 -549
rect 77 -557 81 -552
rect 72 -561 81 -557
rect 48 -576 52 -573
rect 87 -576 91 -541
rect 99 -542 103 -534
rect 28 -582 38 -578
rect 48 -580 91 -576
rect 59 -588 63 -580
rect 37 -603 41 -598
rect 50 -603 52 -599
rect 32 -607 41 -603
rect 30 -614 66 -611
rect 30 -615 56 -614
rect 30 -619 34 -615
rect 52 -619 56 -615
rect 62 -619 66 -614
rect 41 -642 45 -639
rect 74 -642 78 -639
rect 41 -646 65 -642
rect 74 -646 89 -642
rect 29 -648 31 -647
rect -18 -651 31 -648
rect 52 -654 56 -646
rect 74 -654 78 -646
rect 30 -669 34 -664
rect 28 -670 34 -669
rect 62 -670 66 -664
rect 28 -673 66 -670
rect 34 -678 40 -676
rect -27 -681 40 -678
rect 85 -796 89 -646
rect 137 -671 140 -534
rect 144 -543 147 -534
rect 155 -536 159 -531
rect 151 -540 159 -536
rect 162 -543 166 -536
rect 144 -547 166 -543
rect 170 -607 173 -536
rect 185 -571 189 -513
rect 194 -527 198 -522
rect 207 -527 209 -523
rect 223 -525 227 -504
rect 245 -523 249 -520
rect 192 -533 198 -527
rect 223 -529 235 -525
rect 245 -527 262 -523
rect 256 -528 262 -527
rect 244 -534 249 -530
rect 205 -538 209 -535
rect 194 -542 220 -538
rect 194 -546 198 -542
rect 216 -546 220 -542
rect 234 -550 238 -545
rect 229 -554 238 -550
rect 205 -569 209 -566
rect 244 -569 248 -534
rect 256 -535 260 -528
rect 185 -575 195 -571
rect 205 -573 248 -569
rect 216 -581 220 -573
rect 194 -596 198 -591
rect 189 -600 198 -596
rect 209 -598 213 -596
rect 284 -598 287 -459
rect 296 -527 298 -524
rect 209 -601 287 -598
rect 209 -607 212 -601
rect 170 -610 212 -607
rect 359 -621 362 -433
rect 155 -624 362 -621
rect 155 -627 160 -624
rect 207 -631 308 -628
rect 207 -634 211 -631
rect 304 -634 308 -631
rect 146 -638 182 -635
rect 146 -639 172 -638
rect 146 -643 150 -639
rect 168 -643 172 -639
rect 178 -643 182 -638
rect 197 -638 211 -634
rect 219 -638 255 -635
rect 157 -666 161 -663
rect 190 -666 194 -663
rect 197 -664 200 -638
rect 219 -639 245 -638
rect 219 -643 223 -639
rect 241 -643 245 -639
rect 251 -643 255 -638
rect 270 -638 291 -634
rect 157 -670 181 -666
rect 190 -670 197 -666
rect 230 -666 234 -663
rect 263 -666 267 -663
rect 270 -665 273 -638
rect 286 -644 319 -641
rect 286 -645 293 -644
rect 289 -648 293 -645
rect 315 -648 319 -644
rect 230 -670 254 -666
rect 263 -670 270 -666
rect 137 -675 147 -671
rect 137 -704 140 -675
rect 160 -677 161 -673
rect 168 -678 172 -670
rect 190 -678 194 -670
rect 213 -675 220 -671
rect 146 -694 150 -688
rect 178 -694 182 -688
rect 146 -697 182 -694
rect 163 -701 170 -697
rect 213 -704 216 -675
rect 233 -677 234 -673
rect 241 -678 245 -670
rect 263 -678 267 -670
rect 306 -671 310 -668
rect 323 -671 327 -668
rect 298 -675 316 -671
rect 323 -674 334 -671
rect 298 -680 302 -675
rect 323 -680 327 -674
rect 219 -694 223 -688
rect 251 -694 255 -688
rect 219 -697 255 -694
rect 289 -694 293 -690
rect 307 -694 311 -690
rect 315 -694 319 -690
rect 289 -697 319 -694
rect 236 -701 243 -697
rect 302 -700 305 -697
rect 137 -707 216 -704
rect 330 -709 334 -674
rect 244 -712 334 -709
rect 244 -715 248 -712
rect 261 -719 298 -715
rect 239 -725 272 -722
rect 239 -726 246 -725
rect 242 -729 246 -726
rect 268 -729 272 -725
rect 259 -752 263 -749
rect 276 -752 280 -749
rect 251 -756 269 -752
rect 276 -755 284 -752
rect 251 -761 255 -756
rect 276 -761 280 -755
rect 242 -775 246 -771
rect 260 -775 264 -771
rect 268 -775 272 -771
rect 242 -778 272 -775
rect 255 -781 258 -778
rect 295 -796 298 -719
rect 85 -799 352 -796
rect 285 -837 288 -809
rect 284 -840 288 -837
rect 177 -853 238 -849
rect 20 -860 81 -856
rect 177 -858 181 -853
rect 20 -865 24 -860
rect -6 -869 24 -865
rect -2 -873 2 -869
rect 20 -873 24 -869
rect -38 -880 -15 -877
rect -38 -889 -24 -886
rect -27 -936 -24 -889
rect -18 -910 -15 -880
rect 37 -864 41 -860
rect 59 -864 63 -860
rect 77 -879 81 -860
rect 155 -862 181 -858
rect 155 -866 159 -862
rect 177 -866 181 -862
rect 77 -883 103 -879
rect 48 -887 52 -884
rect 77 -887 81 -883
rect 99 -887 103 -883
rect 194 -857 198 -853
rect 216 -857 220 -853
rect 234 -872 238 -853
rect 234 -876 260 -872
rect 205 -880 209 -877
rect 234 -880 238 -876
rect 256 -880 260 -876
rect 205 -884 227 -880
rect 48 -891 70 -887
rect 9 -896 13 -893
rect 28 -895 38 -891
rect 28 -896 32 -895
rect 9 -900 32 -896
rect 59 -899 63 -891
rect 20 -908 24 -900
rect -18 -928 -15 -915
rect -2 -923 2 -918
rect -6 -927 2 -923
rect 5 -930 9 -923
rect -13 -933 9 -930
rect 13 -936 17 -923
rect -27 -939 17 -936
rect -27 -979 -24 -939
rect -27 -1058 -24 -984
rect -18 -1028 -15 -950
rect 28 -958 32 -900
rect 37 -914 41 -909
rect 35 -920 41 -914
rect 66 -912 70 -891
rect 166 -889 170 -886
rect 185 -888 195 -884
rect 185 -889 189 -888
rect 166 -893 189 -889
rect 216 -892 220 -884
rect 177 -901 181 -893
rect 88 -910 92 -907
rect 142 -910 147 -908
rect 66 -916 78 -912
rect 88 -914 147 -910
rect 87 -921 92 -917
rect 48 -925 52 -922
rect 37 -929 63 -925
rect 37 -933 41 -929
rect 59 -933 63 -929
rect 77 -937 81 -932
rect 72 -941 81 -937
rect 48 -956 52 -953
rect 87 -956 91 -921
rect 99 -922 103 -914
rect 28 -962 38 -958
rect 48 -960 91 -956
rect 59 -968 63 -960
rect 37 -983 41 -978
rect 32 -987 41 -983
rect 30 -994 66 -991
rect 30 -995 56 -994
rect 30 -999 34 -995
rect 52 -999 56 -995
rect 62 -999 66 -994
rect 41 -1022 45 -1019
rect 74 -1022 78 -1019
rect 41 -1026 65 -1022
rect 74 -1026 89 -1022
rect 29 -1028 31 -1027
rect -18 -1031 31 -1028
rect 52 -1034 56 -1026
rect 74 -1034 78 -1026
rect 30 -1049 34 -1044
rect 28 -1050 34 -1049
rect 62 -1050 66 -1044
rect 28 -1053 66 -1050
rect 34 -1058 40 -1056
rect -27 -1061 40 -1058
rect 85 -1194 89 -1026
rect 137 -1051 140 -914
rect 144 -923 147 -914
rect 155 -916 159 -911
rect 151 -920 159 -916
rect 162 -923 166 -916
rect 144 -927 166 -923
rect 170 -987 173 -916
rect 185 -951 189 -893
rect 194 -907 198 -902
rect 192 -913 198 -907
rect 223 -905 227 -884
rect 245 -903 249 -900
rect 223 -909 235 -905
rect 245 -907 262 -903
rect 256 -908 262 -907
rect 244 -914 249 -910
rect 205 -918 209 -915
rect 194 -922 220 -918
rect 194 -926 198 -922
rect 216 -926 220 -922
rect 234 -930 238 -925
rect 229 -934 238 -930
rect 205 -949 209 -946
rect 244 -949 248 -914
rect 256 -915 260 -908
rect 185 -955 195 -951
rect 205 -953 248 -949
rect 216 -961 220 -953
rect 194 -976 198 -971
rect 189 -980 198 -976
rect 209 -978 213 -976
rect 284 -978 287 -840
rect 296 -907 298 -904
rect 209 -981 287 -978
rect 209 -987 212 -981
rect 170 -990 212 -987
rect 349 -1001 352 -799
rect 155 -1004 352 -1001
rect 155 -1007 160 -1004
rect 207 -1011 309 -1008
rect 207 -1014 211 -1011
rect 305 -1014 309 -1011
rect 146 -1018 182 -1015
rect 146 -1019 172 -1018
rect 146 -1023 150 -1019
rect 168 -1023 172 -1019
rect 178 -1023 182 -1018
rect 197 -1018 211 -1014
rect 219 -1018 255 -1015
rect 157 -1046 161 -1043
rect 190 -1046 194 -1043
rect 197 -1046 200 -1018
rect 219 -1019 245 -1018
rect 219 -1023 223 -1019
rect 241 -1023 245 -1019
rect 251 -1023 255 -1018
rect 270 -1018 292 -1014
rect 157 -1050 181 -1046
rect 190 -1050 200 -1046
rect 230 -1046 234 -1043
rect 263 -1046 267 -1043
rect 270 -1046 273 -1018
rect 287 -1024 320 -1021
rect 287 -1025 294 -1024
rect 230 -1050 254 -1046
rect 263 -1050 273 -1046
rect 290 -1028 294 -1025
rect 316 -1028 320 -1024
rect 137 -1055 147 -1051
rect 137 -1084 140 -1055
rect 160 -1057 161 -1053
rect 168 -1058 172 -1050
rect 190 -1058 194 -1050
rect 213 -1055 220 -1051
rect 146 -1074 150 -1068
rect 178 -1074 182 -1068
rect 146 -1077 182 -1074
rect 163 -1081 170 -1077
rect 213 -1084 216 -1055
rect 233 -1057 234 -1053
rect 241 -1058 245 -1050
rect 263 -1058 267 -1050
rect 307 -1051 311 -1048
rect 324 -1051 328 -1048
rect 299 -1055 317 -1051
rect 324 -1054 335 -1051
rect 299 -1060 303 -1055
rect 324 -1060 328 -1054
rect 219 -1074 223 -1068
rect 251 -1074 255 -1068
rect 219 -1077 255 -1074
rect 290 -1074 294 -1070
rect 308 -1074 312 -1070
rect 316 -1074 320 -1070
rect 290 -1077 320 -1074
rect 236 -1081 243 -1077
rect 303 -1080 306 -1077
rect 137 -1087 216 -1084
rect 137 -1143 141 -1087
rect 331 -1106 335 -1054
rect 144 -1110 180 -1107
rect 144 -1111 170 -1110
rect 144 -1115 148 -1111
rect 166 -1115 170 -1111
rect 176 -1115 180 -1110
rect 195 -1110 211 -1106
rect 228 -1110 335 -1106
rect 155 -1138 159 -1135
rect 188 -1138 192 -1135
rect 195 -1138 198 -1110
rect 206 -1116 239 -1113
rect 206 -1117 213 -1116
rect 155 -1142 179 -1138
rect 188 -1142 198 -1138
rect 209 -1120 213 -1117
rect 235 -1120 239 -1116
rect 251 -1117 261 -1113
rect 278 -1117 315 -1113
rect 137 -1147 145 -1143
rect 158 -1149 159 -1145
rect 166 -1150 170 -1142
rect 188 -1150 192 -1142
rect 226 -1143 230 -1140
rect 243 -1143 247 -1140
rect 251 -1143 254 -1117
rect 218 -1147 236 -1143
rect 243 -1146 254 -1143
rect 259 -1123 289 -1120
rect 259 -1127 263 -1123
rect 285 -1127 289 -1123
rect 218 -1152 222 -1147
rect 243 -1152 247 -1146
rect 276 -1150 280 -1147
rect 144 -1166 148 -1160
rect 176 -1166 180 -1160
rect 144 -1169 180 -1166
rect 209 -1166 213 -1162
rect 227 -1166 231 -1162
rect 268 -1154 286 -1150
rect 268 -1159 272 -1154
rect 293 -1159 297 -1147
rect 235 -1166 239 -1162
rect 209 -1169 239 -1166
rect 161 -1173 168 -1169
rect 222 -1172 225 -1169
rect 259 -1173 263 -1169
rect 277 -1173 281 -1169
rect 285 -1173 289 -1169
rect 259 -1176 289 -1173
rect 272 -1179 275 -1176
rect 312 -1194 315 -1117
rect 354 -1154 358 -1151
rect 85 -1197 315 -1194
rect 227 -1345 236 -1342
<< m2contact >>
rect 123 40 128 45
rect 123 -6 128 -1
rect -23 -19 -18 -14
rect -23 -36 -18 -31
rect 289 6 294 11
rect 318 6 323 11
rect 35 -120 40 -115
rect 35 -147 40 -142
rect 202 -166 207 -161
rect -24 -268 -19 -263
rect -24 -285 -19 -280
rect 34 -369 39 -364
rect 34 -396 39 -391
rect 256 -243 261 -238
rect 298 -166 303 -161
rect 285 -243 290 -238
rect 149 -347 154 -342
rect 191 -385 196 -380
rect 149 -393 154 -388
rect 255 -390 260 -385
rect 255 -443 260 -438
rect -18 -553 -13 -548
rect -18 -570 -13 -565
rect 40 -654 45 -649
rect 40 -681 45 -676
rect 262 -528 267 -523
rect 291 -528 296 -523
rect 155 -632 160 -627
rect 197 -670 203 -664
rect 270 -670 275 -665
rect 155 -678 160 -673
rect 228 -678 233 -673
rect 284 -756 289 -751
rect 284 -809 289 -804
rect -18 -915 -13 -910
rect -18 -933 -13 -928
rect -29 -984 -24 -979
rect -18 -950 -13 -945
rect 47 -915 52 -910
rect 142 -908 147 -903
rect 47 -984 52 -979
rect 40 -1034 45 -1029
rect 40 -1061 45 -1056
rect 204 -908 209 -903
rect 262 -908 267 -903
rect 291 -908 296 -903
rect 155 -1012 160 -1007
rect 155 -1058 160 -1053
rect 228 -1058 233 -1053
rect 153 -1150 158 -1145
rect 297 -1155 302 -1150
rect 349 -1155 354 -1150
<< metal2 >>
rect 123 -1 128 40
rect 294 7 318 10
rect -23 -31 -18 -19
rect 35 -142 40 -120
rect 207 -166 298 -161
rect 261 -242 285 -239
rect -24 -280 -19 -268
rect 34 -391 39 -369
rect 149 -388 154 -347
rect 191 -453 196 -385
rect 255 -438 260 -390
rect 191 -456 233 -453
rect -18 -565 -13 -553
rect 40 -676 45 -654
rect 155 -673 160 -632
rect 198 -838 201 -670
rect 228 -673 233 -456
rect 267 -527 291 -524
rect 198 -842 233 -838
rect 147 -907 155 -904
rect 202 -907 204 -904
rect -13 -914 47 -911
rect -18 -945 -13 -933
rect -24 -983 47 -980
rect 40 -1056 45 -1034
rect 155 -1053 160 -1012
rect 228 -1053 233 -842
rect 271 -894 274 -670
rect 284 -804 289 -756
rect 271 -897 303 -894
rect 267 -907 291 -904
rect 300 -931 303 -897
rect 250 -934 303 -931
rect 250 -1101 253 -934
rect 153 -1104 253 -1101
rect 153 -1145 158 -1104
rect 302 -1154 349 -1151
use xor  xor_0
timestamp 1618484725
transform 1 0 0 0 1 -22
box -11 -51 105 80
use and  and_1
timestamp 1618590203
transform 1 0 111 0 1 -25
box 1 0 54 62
use xor  xor_1
timestamp 1618484725
transform 1 0 189 0 1 -15
box -11 -51 105 80
use and  and_0
timestamp 1618590203
transform 1 0 22 0 1 -139
box 1 0 54 62
use or  or_0
timestamp 1618732609
transform 1 0 118 0 1 -112
box -27 -27 14 35
<< labels >>
rlabel metal1 -39 35 -39 35 3 a1
rlabel metal1 -38 26 -38 26 3 b1
rlabel metal1 46 2 46 2 1 a1
rlabel metal1 46 -67 46 -67 1 b1
rlabel metal1 110 1 110 1 1 p1
rlabel metal1 166 4 166 4 1 i1
rlabel metal1 77 -110 77 -110 1 g1
rlabel metal1 235 9 235 9 1 p1
rlabel metal1 325 9 325 9 7 sum1
rlabel metal1 125 46 125 46 1 c0
rlabel metal1 312 75 312 75 5 c0
rlabel metal1 -40 -213 -40 -213 3 a2
rlabel metal1 -37 -222 -37 -222 1 b2
rlabel metal1 42 -194 42 -194 1 vdd
rlabel metal1 45 -262 45 -262 1 vdd
rlabel metal1 34 -250 34 -250 1 gnd
rlabel metal1 -8 -261 -8 -261 1 gnd
rlabel metal1 70 -274 70 -274 1 gnd
rlabel metal1 33 -318 33 -318 1 gnd
rlabel metal1 25 -385 25 -385 1 gnd
rlabel metal1 37 -328 37 -328 1 vdd
rlabel metal1 45 -247 45 -247 1 a2
rlabel metal1 45 -316 45 -316 1 b2
rlabel metal1 99 -248 99 -248 1 p2
rlabel metal1 74 -359 74 -359 1 g2
rlabel metal1 41 61 41 61 1 vdd
rlabel metal1 51 -10 51 -10 1 vdd
rlabel metal1 46 -76 46 -76 1 vdd
rlabel metal1 113 36 113 36 1 vdd
rlabel metal1 231 66 231 66 1 vdd
rlabel metal1 239 -2 239 -2 1 vdd
rlabel metal1 34 -7 34 -7 1 gnd
rlabel metal1 72 -28 72 -28 1 gnd
rlabel metal1 -12 -10 -12 -10 1 gnd
rlabel metal1 54 -140 54 -140 1 gnd
rlabel metal1 106 -140 106 -140 1 gnd
rlabel metal1 136 -28 136 -28 1 gnd
rlabel metal1 180 -1 180 -1 1 gnd
rlabel metal1 90 -85 90 -85 1 vdd
rlabel metal1 226 3 226 3 1 gnd
rlabel metal1 260 -21 260 -21 1 gnd
rlabel metal1 215 -64 215 -64 1 gnd
rlabel metal1 205 -186 205 -186 1 vdd
rlabel metal1 202 -253 202 -253 1 vdd
rlabel metal1 189 -313 189 -313 1 gnd
rlabel metal1 149 -253 149 -253 1 gnd
rlabel metal1 191 -246 191 -246 1 gnd
rlabel metal1 229 -268 229 -268 1 gnd
rlabel metal1 291 -240 291 -240 7 sum2
rlabel metal1 202 -240 202 -240 1 p2
rlabel metal1 142 -351 142 -351 1 vdd
rlabel metal1 160 -414 160 -414 1 gnd
rlabel metal1 228 -414 228 -414 1 gnd
rlabel metal1 236 -358 236 -358 1 vdd
rlabel metal1 253 -387 253 -387 1 c2
rlabel metal1 48 -479 48 -479 1 vdd
rlabel metal1 51 -547 51 -547 1 vdd
rlabel metal1 40 -535 40 -535 1 gnd
rlabel metal1 -2 -546 -2 -546 1 gnd
rlabel metal1 76 -559 76 -559 1 gnd
rlabel metal1 39 -603 39 -603 1 gnd
rlabel metal1 31 -670 31 -670 1 gnd
rlabel metal1 43 -613 43 -613 1 vdd
rlabel metal1 211 -471 211 -471 1 vdd
rlabel metal1 208 -538 208 -538 1 vdd
rlabel metal1 195 -598 195 -598 1 gnd
rlabel metal1 155 -538 155 -538 1 gnd
rlabel metal1 197 -531 197 -531 1 gnd
rlabel metal1 235 -553 235 -553 1 gnd
rlabel metal1 148 -636 148 -636 1 vdd
rlabel metal1 166 -699 166 -699 1 gnd
rlabel metal1 -30 -499 -30 -499 1 a3
rlabel metal1 -32 -508 -32 -508 1 b3
rlabel metal1 51 -532 51 -532 1 a3
rlabel metal1 51 -602 51 -602 1 b3
rlabel metal1 113 -532 113 -532 1 p3
rlabel metal1 297 -526 297 -526 1 sum3
rlabel metal1 136 -114 136 -114 1 c1
rlabel metal1 239 -699 239 -699 1 gnd
rlabel metal1 221 -636 221 -636 1 vdd
rlabel metal1 304 -699 304 -699 1 gnd
rlabel metal1 312 -643 312 -643 1 vdd
rlabel metal1 257 -780 257 -780 1 gnd
rlabel metal1 265 -724 265 -724 1 vdd
rlabel metal1 282 -754 282 -754 1 c3
rlabel metal1 208 -524 208 -524 1 p3
rlabel metal1 48 -859 48 -859 1 vdd
rlabel metal1 51 -927 51 -927 1 vdd
rlabel metal1 40 -915 40 -915 1 gnd
rlabel metal1 -2 -926 -2 -926 1 gnd
rlabel metal1 76 -939 76 -939 1 gnd
rlabel metal1 39 -983 39 -983 1 gnd
rlabel metal1 31 -1050 31 -1050 1 gnd
rlabel metal1 43 -993 43 -993 1 vdd
rlabel metal1 211 -851 211 -851 1 vdd
rlabel metal1 208 -918 208 -918 1 vdd
rlabel metal1 195 -978 195 -978 1 gnd
rlabel metal1 155 -918 155 -918 1 gnd
rlabel metal1 197 -911 197 -911 1 gnd
rlabel metal1 235 -933 235 -933 1 gnd
rlabel metal1 148 -1016 148 -1016 1 vdd
rlabel metal1 166 -1079 166 -1079 1 gnd
rlabel metal1 239 -1079 239 -1079 1 gnd
rlabel metal1 221 -1016 221 -1016 1 vdd
rlabel metal1 -33 -878 -33 -878 1 a4
rlabel metal1 -33 -887 -33 -887 1 b4
rlabel metal1 116 -913 116 -913 1 p4
rlabel metal1 82 -1025 82 -1025 1 g4
rlabel metal1 81 -645 81 -645 1 g3
rlabel metal1 146 -1108 146 -1108 1 vdd
rlabel metal1 164 -1171 164 -1171 1 gnd
rlabel metal1 305 -1079 305 -1079 1 gnd
rlabel metal1 313 -1023 313 -1023 1 vdd
rlabel metal1 224 -1171 224 -1171 1 gnd
rlabel metal1 232 -1115 232 -1115 1 vdd
rlabel metal1 274 -1178 274 -1178 1 gnd
rlabel metal1 282 -1122 282 -1122 1 vdd
rlabel metal1 356 -1153 356 -1153 1 cout
rlabel metal1 297 -906 297 -906 1 sum4
rlabel metal2 203 -906 203 -906 1 p4
<< end >>
